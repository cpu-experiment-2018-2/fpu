`default_nettype none

module fdiv(
input wire [31:0] adata,
input wire [31:0] bdata,
output reg [31:0] result,
input wire clk,
input wire flag_in,
input wire [4:0] address_in,
output reg flag_out,
output reg [4:0] address_out);

(* ram_style = "distributed" *) reg [22:0] key [1024:0];
(* ram_style = "distributed" *) reg [12:0] key2 [1024:0];
(* ram_style = "distributed" *) reg key3 [1024:0];


assign key[0] = 8388607;
assign key2[0] = 8190;
assign key3[0] = 0;
assign key[1] = 8372242;
assign key2[1] = 8176;
assign key3[1] = 0;
assign key[2] = 8355906;
assign key2[2] = 8160;
assign key3[2] = 0;
assign key[3] = 8339602;
assign key2[3] = 8144;
assign key3[3] = 0;
assign key[4] = 8323329;
assign key2[4] = 8128;
assign key3[4] = 0;
assign key[5] = 8307088;
assign key2[5] = 8112;
assign key3[5] = 0;
assign key[6] = 8290879;
assign key2[6] = 8096;
assign key3[6] = 0;
assign key[7] = 8274701;
assign key2[7] = 8081;
assign key3[7] = 0;
assign key[8] = 8258554;
assign key2[8] = 8065;
assign key3[8] = 0;
assign key[9] = 8242439;
assign key2[9] = 8049;
assign key3[9] = 0;
assign key[10] = 8226354;
assign key2[10] = 8034;
assign key3[10] = 0;
assign key[11] = 8210301;
assign key2[11] = 8018;
assign key3[11] = 0;
assign key[12] = 8194279;
assign key2[12] = 8003;
assign key3[12] = 0;
assign key[13] = 8178288;
assign key2[13] = 7987;
assign key3[13] = 0;
assign key[14] = 8162328;
assign key2[14] = 7972;
assign key3[14] = 0;
assign key[15] = 8146398;
assign key2[15] = 7957;
assign key3[15] = 0;
assign key[16] = 8130499;
assign key2[16] = 7941;
assign key3[16] = 0;
assign key[17] = 8114630;
assign key2[17] = 7926;
assign key3[17] = 0;
assign key[18] = 8098792;
assign key2[18] = 7911;
assign key3[18] = 0;
assign key[19] = 8082985;
assign key2[19] = 7896;
assign key3[19] = 0;
assign key[20] = 8067207;
assign key2[20] = 7881;
assign key3[20] = 0;
assign key[21] = 8051460;
assign key2[21] = 7866;
assign key3[21] = 0;
assign key[22] = 8035743;
assign key2[22] = 7851;
assign key3[22] = 0;
assign key[23] = 8020056;
assign key2[23] = 7836;
assign key3[23] = 0;
assign key[24] = 8004399;
assign key2[24] = 7821;
assign key3[24] = 0;
assign key[25] = 7988772;
assign key2[25] = 7806;
assign key3[25] = 0;
assign key[26] = 7973174;
assign key2[26] = 7791;
assign key3[26] = 0;
assign key[27] = 7957606;
assign key2[27] = 7776;
assign key3[27] = 0;
assign key[28] = 7942068;
assign key2[28] = 7761;
assign key3[28] = 0;
assign key[29] = 7926559;
assign key2[29] = 7746;
assign key3[29] = 0;
assign key[30] = 7911080;
assign key2[30] = 7732;
assign key3[30] = 0;
assign key[31] = 7895630;
assign key2[31] = 7717;
assign key3[31] = 0;
assign key[32] = 7880209;
assign key2[32] = 7703;
assign key3[32] = 0;
assign key[33] = 7864818;
assign key2[33] = 7688;
assign key3[33] = 0;
assign key[34] = 7849455;
assign key2[34] = 7673;
assign key3[34] = 0;
assign key[35] = 7834122;
assign key2[35] = 7659;
assign key3[35] = 0;
assign key[36] = 7818818;
assign key2[36] = 7645;
assign key3[36] = 0;
assign key[37] = 7803542;
assign key2[37] = 7630;
assign key3[37] = 0;
assign key[38] = 7788295;
assign key2[38] = 7616;
assign key3[38] = 0;
assign key[39] = 7773077;
assign key2[39] = 7601;
assign key3[39] = 0;
assign key[40] = 7757887;
assign key2[40] = 7587;
assign key3[40] = 0;
assign key[41] = 7742726;
assign key2[41] = 7573;
assign key3[41] = 0;
assign key[42] = 7727594;
assign key2[42] = 7559;
assign key3[42] = 0;
assign key[43] = 7712490;
assign key2[43] = 7545;
assign key3[43] = 0;
assign key[44] = 7697414;
assign key2[44] = 7530;
assign key3[44] = 0;
assign key[45] = 7682366;
assign key2[45] = 7516;
assign key3[45] = 0;
assign key[46] = 7667346;
assign key2[46] = 7502;
assign key3[46] = 0;
assign key[47] = 7652355;
assign key2[47] = 7488;
assign key3[47] = 0;
assign key[48] = 7637391;
assign key2[48] = 7474;
assign key3[48] = 0;
assign key[49] = 7622455;
assign key2[49] = 7460;
assign key3[49] = 0;
assign key[50] = 7607548;
assign key2[50] = 7446;
assign key3[50] = 0;
assign key[51] = 7592667;
assign key2[51] = 7433;
assign key3[51] = 0;
assign key[52] = 7577815;
assign key2[52] = 7419;
assign key3[52] = 0;
assign key[53] = 7562990;
assign key2[53] = 7405;
assign key3[53] = 0;
assign key[54] = 7548193;
assign key2[54] = 7391;
assign key3[54] = 0;
assign key[55] = 7533423;
assign key2[55] = 7378;
assign key3[55] = 0;
assign key[56] = 7518680;
assign key2[56] = 7364;
assign key3[56] = 0;
assign key[57] = 7503965;
assign key2[57] = 7350;
assign key3[57] = 0;
assign key[58] = 7489276;
assign key2[58] = 7337;
assign key3[58] = 0;
assign key[59] = 7474615;
assign key2[59] = 7323;
assign key3[59] = 0;
assign key[60] = 7459981;
assign key2[60] = 7310;
assign key3[60] = 0;
assign key[61] = 7445374;
assign key2[61] = 7296;
assign key3[61] = 0;
assign key[62] = 7430794;
assign key2[62] = 7283;
assign key3[62] = 0;
assign key[63] = 7416241;
assign key2[63] = 7269;
assign key3[63] = 0;
assign key[64] = 7401715;
assign key2[64] = 7256;
assign key3[64] = 0;
assign key[65] = 7387215;
assign key2[65] = 7243;
assign key3[65] = 0;
assign key[66] = 7372742;
assign key2[66] = 7229;
assign key3[66] = 0;
assign key[67] = 7358295;
assign key2[67] = 7216;
assign key3[67] = 0;
assign key[68] = 7343875;
assign key2[68] = 7203;
assign key3[68] = 0;
assign key[69] = 7329481;
assign key2[69] = 7190;
assign key3[69] = 0;
assign key[70] = 7315113;
assign key2[70] = 7177;
assign key3[70] = 0;
assign key[71] = 7300772;
assign key2[71] = 7164;
assign key3[71] = 0;
assign key[72] = 7286457;
assign key2[72] = 7151;
assign key3[72] = 0;
assign key[73] = 7272168;
assign key2[73] = 7138;
assign key3[73] = 0;
assign key[74] = 7257905;
assign key2[74] = 7125;
assign key3[74] = 0;
assign key[75] = 7243668;
assign key2[75] = 7112;
assign key3[75] = 0;
assign key[76] = 7229457;
assign key2[76] = 7099;
assign key3[76] = 0;
assign key[77] = 7215271;
assign key2[77] = 7086;
assign key3[77] = 0;
assign key[78] = 7201112;
assign key2[78] = 7073;
assign key3[78] = 0;
assign key[79] = 7186978;
assign key2[79] = 7060;
assign key3[79] = 0;
assign key[80] = 7172869;
assign key2[80] = 7047;
assign key3[80] = 0;
assign key[81] = 7158787;
assign key2[81] = 7035;
assign key3[81] = 0;
assign key[82] = 7144729;
assign key2[82] = 7022;
assign key3[82] = 0;
assign key[83] = 7130697;
assign key2[83] = 7009;
assign key3[83] = 0;
assign key[84] = 7116691;
assign key2[84] = 6996;
assign key3[84] = 0;
assign key[85] = 7102709;
assign key2[85] = 6984;
assign key3[85] = 0;
assign key[86] = 7088753;
assign key2[86] = 6971;
assign key3[86] = 0;
assign key[87] = 7074822;
assign key2[87] = 6959;
assign key3[87] = 0;
assign key[88] = 7060916;
assign key2[88] = 6946;
assign key3[88] = 0;
assign key[89] = 7047035;
assign key2[89] = 6934;
assign key3[89] = 0;
assign key[90] = 7033179;
assign key2[90] = 6921;
assign key3[90] = 0;
assign key[91] = 7019348;
assign key2[91] = 6909;
assign key3[91] = 0;
assign key[92] = 7005542;
assign key2[92] = 6897;
assign key3[92] = 0;
assign key[93] = 6991760;
assign key2[93] = 6884;
assign key3[93] = 0;
assign key[94] = 6978003;
assign key2[94] = 6872;
assign key3[94] = 0;
assign key[95] = 6964270;
assign key2[95] = 6860;
assign key3[95] = 0;
assign key[96] = 6950562;
assign key2[96] = 6847;
assign key3[96] = 0;
assign key[97] = 6936879;
assign key2[97] = 6835;
assign key3[97] = 0;
assign key[98] = 6923220;
assign key2[98] = 6823;
assign key3[98] = 0;
assign key[99] = 6909585;
assign key2[99] = 6811;
assign key3[99] = 0;
assign key[100] = 6895975;
assign key2[100] = 6799;
assign key3[100] = 0;
assign key[101] = 6882388;
assign key2[101] = 6787;
assign key3[101] = 0;
assign key[102] = 6868826;
assign key2[102] = 6775;
assign key3[102] = 0;
assign key[103] = 6855288;
assign key2[103] = 6763;
assign key3[103] = 0;
assign key[104] = 6841774;
assign key2[104] = 6751;
assign key3[104] = 0;
assign key[105] = 6828284;
assign key2[105] = 6739;
assign key3[105] = 0;
assign key[106] = 6814818;
assign key2[106] = 6727;
assign key3[106] = 0;
assign key[107] = 6801375;
assign key2[107] = 6715;
assign key3[107] = 0;
assign key[108] = 6787956;
assign key2[108] = 6703;
assign key3[108] = 0;
assign key[109] = 6774561;
assign key2[109] = 6691;
assign key3[109] = 0;
assign key[110] = 6761190;
assign key2[110] = 6679;
assign key3[110] = 0;
assign key[111] = 6747842;
assign key2[111] = 6668;
assign key3[111] = 0;
assign key[112] = 6734518;
assign key2[112] = 6656;
assign key3[112] = 0;
assign key[113] = 6721217;
assign key2[113] = 6644;
assign key3[113] = 0;
assign key[114] = 6707939;
assign key2[114] = 6632;
assign key3[114] = 0;
assign key[115] = 6694685;
assign key2[115] = 6621;
assign key3[115] = 0;
assign key[116] = 6681454;
assign key2[116] = 6609;
assign key3[116] = 0;
assign key[117] = 6668246;
assign key2[117] = 6598;
assign key3[117] = 0;
assign key[118] = 6655062;
assign key2[118] = 6586;
assign key3[118] = 0;
assign key[119] = 6641900;
assign key2[119] = 6575;
assign key3[119] = 0;
assign key[120] = 6628762;
assign key2[120] = 6563;
assign key3[120] = 0;
assign key[121] = 6615646;
assign key2[121] = 6552;
assign key3[121] = 0;
assign key[122] = 6602553;
assign key2[122] = 6540;
assign key3[122] = 0;
assign key[123] = 6589483;
assign key2[123] = 6529;
assign key3[123] = 0;
assign key[124] = 6576436;
assign key2[124] = 6517;
assign key3[124] = 0;
assign key[125] = 6563412;
assign key2[125] = 6506;
assign key3[125] = 0;
assign key[126] = 6550410;
assign key2[126] = 6495;
assign key3[126] = 0;
assign key[127] = 6537431;
assign key2[127] = 6483;
assign key3[127] = 0;
assign key[128] = 6524474;
assign key2[128] = 6472;
assign key3[128] = 0;
assign key[129] = 6511540;
assign key2[129] = 6461;
assign key3[129] = 0;
assign key[130] = 6498628;
assign key2[130] = 6450;
assign key3[130] = 0;
assign key[131] = 6485739;
assign key2[131] = 6439;
assign key3[131] = 0;
assign key[132] = 6472872;
assign key2[132] = 6427;
assign key3[132] = 0;
assign key[133] = 6460027;
assign key2[133] = 6416;
assign key3[133] = 0;
assign key[134] = 6447204;
assign key2[134] = 6405;
assign key3[134] = 0;
assign key[135] = 6434404;
assign key2[135] = 6394;
assign key3[135] = 0;
assign key[136] = 6421625;
assign key2[136] = 6383;
assign key3[136] = 0;
assign key[137] = 6408869;
assign key2[137] = 6372;
assign key3[137] = 0;
assign key[138] = 6396134;
assign key2[138] = 6361;
assign key3[138] = 0;
assign key[139] = 6383422;
assign key2[139] = 6350;
assign key3[139] = 0;
assign key[140] = 6370731;
assign key2[140] = 6339;
assign key3[140] = 0;
assign key[141] = 6358062;
assign key2[141] = 6329;
assign key3[141] = 0;
assign key[142] = 6345415;
assign key2[142] = 6318;
assign key3[142] = 0;
assign key[143] = 6332789;
assign key2[143] = 6307;
assign key3[143] = 0;
assign key[144] = 6320185;
assign key2[144] = 6296;
assign key3[144] = 0;
assign key[145] = 6307603;
assign key2[145] = 6285;
assign key3[145] = 0;
assign key[146] = 6295042;
assign key2[146] = 6275;
assign key3[146] = 0;
assign key[147] = 6282503;
assign key2[147] = 6264;
assign key3[147] = 0;
assign key[148] = 6269985;
assign key2[148] = 6253;
assign key3[148] = 0;
assign key[149] = 6257488;
assign key2[149] = 6243;
assign key3[149] = 0;
assign key[150] = 6245013;
assign key2[150] = 6232;
assign key3[150] = 0;
assign key[151] = 6232559;
assign key2[151] = 6221;
assign key3[151] = 0;
assign key[152] = 6220126;
assign key2[152] = 6211;
assign key3[152] = 0;
assign key[153] = 6207714;
assign key2[153] = 6200;
assign key3[153] = 0;
assign key[154] = 6195323;
assign key2[154] = 6190;
assign key3[154] = 0;
assign key[155] = 6182953;
assign key2[155] = 6179;
assign key3[155] = 0;
assign key[156] = 6170604;
assign key2[156] = 6169;
assign key3[156] = 0;
assign key[157] = 6158277;
assign key2[157] = 6158;
assign key3[157] = 0;
assign key[158] = 6145970;
assign key2[158] = 6148;
assign key3[158] = 0;
assign key[159] = 6133683;
assign key2[159] = 6137;
assign key3[159] = 0;
assign key[160] = 6121418;
assign key2[160] = 6127;
assign key3[160] = 0;
assign key[161] = 6109173;
assign key2[161] = 6117;
assign key3[161] = 0;
assign key[162] = 6096949;
assign key2[162] = 6106;
assign key3[162] = 0;
assign key[163] = 6084746;
assign key2[163] = 6096;
assign key3[163] = 0;
assign key[164] = 6072563;
assign key2[164] = 6086;
assign key3[164] = 0;
assign key[165] = 6060400;
assign key2[165] = 6076;
assign key3[165] = 0;
assign key[166] = 6048258;
assign key2[166] = 6065;
assign key3[166] = 0;
assign key[167] = 6036136;
assign key2[167] = 6055;
assign key3[167] = 0;
assign key[168] = 6024035;
assign key2[168] = 6045;
assign key3[168] = 0;
assign key[169] = 6011954;
assign key2[169] = 6035;
assign key3[169] = 0;
assign key[170] = 5999893;
assign key2[170] = 6025;
assign key3[170] = 0;
assign key[171] = 5987853;
assign key2[171] = 6015;
assign key3[171] = 0;
assign key[172] = 5975832;
assign key2[172] = 6005;
assign key3[172] = 0;
assign key[173] = 5963832;
assign key2[173] = 5995;
assign key3[173] = 0;
assign key[174] = 5951852;
assign key2[174] = 5985;
assign key3[174] = 0;
assign key[175] = 5939891;
assign key2[175] = 5975;
assign key3[175] = 0;
assign key[176] = 5927951;
assign key2[176] = 5965;
assign key3[176] = 0;
assign key[177] = 5916030;
assign key2[177] = 5955;
assign key3[177] = 0;
assign key[178] = 5904130;
assign key2[178] = 5945;
assign key3[178] = 0;
assign key[179] = 5892249;
assign key2[179] = 5935;
assign key3[179] = 0;
assign key[180] = 5880388;
assign key2[180] = 5925;
assign key3[180] = 0;
assign key[181] = 5868546;
assign key2[181] = 5915;
assign key3[181] = 0;
assign key[182] = 5856724;
assign key2[182] = 5906;
assign key3[182] = 0;
assign key[183] = 5844922;
assign key2[183] = 5896;
assign key3[183] = 0;
assign key[184] = 5833139;
assign key2[184] = 5886;
assign key3[184] = 0;
assign key[185] = 5821376;
assign key2[185] = 5876;
assign key3[185] = 0;
assign key[186] = 5809632;
assign key2[186] = 5867;
assign key3[186] = 0;
assign key[187] = 5797908;
assign key2[187] = 5857;
assign key3[187] = 0;
assign key[188] = 5786203;
assign key2[188] = 5847;
assign key3[188] = 0;
assign key[189] = 5774517;
assign key2[189] = 5838;
assign key3[189] = 0;
assign key[190] = 5762851;
assign key2[190] = 5828;
assign key3[190] = 0;
assign key[191] = 5751203;
assign key2[191] = 5818;
assign key3[191] = 0;
assign key[192] = 5739575;
assign key2[192] = 5809;
assign key3[192] = 0;
assign key[193] = 5727966;
assign key2[193] = 5799;
assign key3[193] = 0;
assign key[194] = 5716376;
assign key2[194] = 5790;
assign key3[194] = 0;
assign key[195] = 5704805;
assign key2[195] = 5780;
assign key3[195] = 0;
assign key[196] = 5693253;
assign key2[196] = 5771;
assign key3[196] = 0;
assign key[197] = 5681720;
assign key2[197] = 5761;
assign key3[197] = 0;
assign key[198] = 5670206;
assign key2[198] = 5752;
assign key3[198] = 0;
assign key[199] = 5658711;
assign key2[199] = 5742;
assign key3[199] = 0;
assign key[200] = 5647234;
assign key2[200] = 5733;
assign key3[200] = 0;
assign key[201] = 5635776;
assign key2[201] = 5724;
assign key3[201] = 0;
assign key[202] = 5624337;
assign key2[202] = 5714;
assign key3[202] = 0;
assign key[203] = 5612917;
assign key2[203] = 5705;
assign key3[203] = 0;
assign key[204] = 5601515;
assign key2[204] = 5696;
assign key3[204] = 0;
assign key[205] = 5590131;
assign key2[205] = 5687;
assign key3[205] = 0;
assign key[206] = 5578766;
assign key2[206] = 5677;
assign key3[206] = 0;
assign key[207] = 5567420;
assign key2[207] = 5668;
assign key3[207] = 0;
assign key[208] = 5556092;
assign key2[208] = 5659;
assign key3[208] = 0;
assign key[209] = 5544783;
assign key2[209] = 5650;
assign key3[209] = 0;
assign key[210] = 5533491;
assign key2[210] = 5641;
assign key3[210] = 0;
assign key[211] = 5522218;
assign key2[211] = 5631;
assign key3[211] = 0;
assign key[212] = 5510964;
assign key2[212] = 5622;
assign key3[212] = 0;
assign key[213] = 5499727;
assign key2[213] = 5613;
assign key3[213] = 0;
assign key[214] = 5488509;
assign key2[214] = 5604;
assign key3[214] = 0;
assign key[215] = 5477309;
assign key2[215] = 5595;
assign key3[215] = 0;
assign key[216] = 5466126;
assign key2[216] = 5586;
assign key3[216] = 0;
assign key[217] = 5454962;
assign key2[217] = 5577;
assign key3[217] = 0;
assign key[218] = 5443816;
assign key2[218] = 5568;
assign key3[218] = 0;
assign key[219] = 5432688;
assign key2[219] = 5559;
assign key3[219] = 0;
assign key[220] = 5421577;
assign key2[220] = 5550;
assign key3[220] = 0;
assign key[221] = 5410485;
assign key2[221] = 5541;
assign key3[221] = 0;
assign key[222] = 5399410;
assign key2[222] = 5532;
assign key3[222] = 0;
assign key[223] = 5388353;
assign key2[223] = 5524;
assign key3[223] = 0;
assign key[224] = 5377314;
assign key2[224] = 5515;
assign key3[224] = 0;
assign key[225] = 5366292;
assign key2[225] = 5506;
assign key3[225] = 0;
assign key[226] = 5355288;
assign key2[226] = 5497;
assign key3[226] = 0;
assign key[227] = 5344302;
assign key2[227] = 5488;
assign key3[227] = 0;
assign key[228] = 5333333;
assign key2[228] = 5480;
assign key3[228] = 0;
assign key[229] = 5322382;
assign key2[229] = 5471;
assign key3[229] = 0;
assign key[230] = 5311448;
assign key2[230] = 5462;
assign key3[230] = 0;
assign key[231] = 5300532;
assign key2[231] = 5453;
assign key3[231] = 0;
assign key[232] = 5289633;
assign key2[232] = 5445;
assign key3[232] = 0;
assign key[233] = 5278751;
assign key2[233] = 5436;
assign key3[233] = 0;
assign key[234] = 5267887;
assign key2[234] = 5427;
assign key3[234] = 0;
assign key[235] = 5257040;
assign key2[235] = 5419;
assign key3[235] = 0;
assign key[236] = 5246210;
assign key2[236] = 5410;
assign key3[236] = 0;
assign key[237] = 5235397;
assign key2[237] = 5402;
assign key3[237] = 0;
assign key[238] = 5224602;
assign key2[238] = 5393;
assign key3[238] = 0;
assign key[239] = 5213823;
assign key2[239] = 5384;
assign key3[239] = 0;
assign key[240] = 5203062;
assign key2[240] = 5376;
assign key3[240] = 0;
assign key[241] = 5192317;
assign key2[241] = 5367;
assign key3[241] = 0;
assign key[242] = 5181590;
assign key2[242] = 5359;
assign key3[242] = 0;
assign key[243] = 5170879;
assign key2[243] = 5351;
assign key3[243] = 0;
assign key[244] = 5160186;
assign key2[244] = 5342;
assign key3[244] = 0;
assign key[245] = 5149509;
assign key2[245] = 5334;
assign key3[245] = 0;
assign key[246] = 5138849;
assign key2[246] = 5325;
assign key3[246] = 0;
assign key[247] = 5128206;
assign key2[247] = 5317;
assign key3[247] = 0;
assign key[248] = 5117580;
assign key2[248] = 5309;
assign key3[248] = 0;
assign key[249] = 5106970;
assign key2[249] = 5300;
assign key3[249] = 0;
assign key[250] = 5096377;
assign key2[250] = 5292;
assign key3[250] = 0;
assign key[251] = 5085800;
assign key2[251] = 5284;
assign key3[251] = 0;
assign key[252] = 5075240;
assign key2[252] = 5275;
assign key3[252] = 0;
assign key[253] = 5064697;
assign key2[253] = 5267;
assign key3[253] = 0;
assign key[254] = 5054170;
assign key2[254] = 5259;
assign key3[254] = 0;
assign key[255] = 5043660;
assign key2[255] = 5251;
assign key3[255] = 0;
assign key[256] = 5033166;
assign key2[256] = 5242;
assign key3[256] = 0;
assign key[257] = 5022688;
assign key2[257] = 5234;
assign key3[257] = 0;
assign key[258] = 5012227;
assign key2[258] = 5226;
assign key3[258] = 0;
assign key[259] = 5001782;
assign key2[259] = 5218;
assign key3[259] = 0;
assign key[260] = 4991353;
assign key2[260] = 5210;
assign key3[260] = 0;
assign key[261] = 4980941;
assign key2[261] = 5202;
assign key3[261] = 0;
assign key[262] = 4970545;
assign key2[262] = 5194;
assign key3[262] = 0;
assign key[263] = 4960165;
assign key2[263] = 5186;
assign key3[263] = 0;
assign key[264] = 4949801;
assign key2[264] = 5177;
assign key3[264] = 0;
assign key[265] = 4939453;
assign key2[265] = 5169;
assign key3[265] = 0;
assign key[266] = 4929121;
assign key2[266] = 5161;
assign key3[266] = 0;
assign key[267] = 4918805;
assign key2[267] = 5153;
assign key3[267] = 0;
assign key[268] = 4908505;
assign key2[268] = 5145;
assign key3[268] = 0;
assign key[269] = 4898221;
assign key2[269] = 5137;
assign key3[269] = 0;
assign key[270] = 4887953;
assign key2[270] = 5130;
assign key3[270] = 0;
assign key[271] = 4877701;
assign key2[271] = 5122;
assign key3[271] = 0;
assign key[272] = 4867465;
assign key2[272] = 5114;
assign key3[272] = 0;
assign key[273] = 4857244;
assign key2[273] = 5106;
assign key3[273] = 0;
assign key[274] = 4847040;
assign key2[274] = 5098;
assign key3[274] = 0;
assign key[275] = 4836850;
assign key2[275] = 5090;
assign key3[275] = 0;
assign key[276] = 4826677;
assign key2[276] = 5082;
assign key3[276] = 0;
assign key[277] = 4816519;
assign key2[277] = 5074;
assign key3[277] = 0;
assign key[278] = 4806377;
assign key2[278] = 5067;
assign key3[278] = 0;
assign key[279] = 4796250;
assign key2[279] = 5059;
assign key3[279] = 0;
assign key[280] = 4786139;
assign key2[280] = 5051;
assign key3[280] = 0;
assign key[281] = 4776044;
assign key2[281] = 5043;
assign key3[281] = 0;
assign key[282] = 4765964;
assign key2[282] = 5036;
assign key3[282] = 0;
assign key[283] = 4755899;
assign key2[283] = 5028;
assign key3[283] = 0;
assign key[284] = 4745850;
assign key2[284] = 5020;
assign key3[284] = 0;
assign key[285] = 4735816;
assign key2[285] = 5013;
assign key3[285] = 0;
assign key[286] = 4725797;
assign key2[286] = 5005;
assign key3[286] = 0;
assign key[287] = 4715794;
assign key2[287] = 4997;
assign key3[287] = 0;
assign key[288] = 4705805;
assign key2[288] = 4990;
assign key3[288] = 0;
assign key[289] = 4695833;
assign key2[289] = 4982;
assign key3[289] = 0;
assign key[290] = 4685875;
assign key2[290] = 4975;
assign key3[290] = 0;
assign key[291] = 4675932;
assign key2[291] = 4967;
assign key3[291] = 0;
assign key[292] = 4666005;
assign key2[292] = 4959;
assign key3[292] = 0;
assign key[293] = 4656092;
assign key2[293] = 4952;
assign key3[293] = 0;
assign key[294] = 4646195;
assign key2[294] = 4944;
assign key3[294] = 0;
assign key[295] = 4636313;
assign key2[295] = 4937;
assign key3[295] = 0;
assign key[296] = 4626445;
assign key2[296] = 4929;
assign key3[296] = 0;
assign key[297] = 4616593;
assign key2[297] = 4922;
assign key3[297] = 0;
assign key[298] = 4606755;
assign key2[298] = 4915;
assign key3[298] = 0;
assign key[299] = 4596933;
assign key2[299] = 4907;
assign key3[299] = 0;
assign key[300] = 4587125;
assign key2[300] = 4900;
assign key3[300] = 0;
assign key[301] = 4577332;
assign key2[301] = 4892;
assign key3[301] = 0;
assign key[302] = 4567554;
assign key2[302] = 4885;
assign key3[302] = 0;
assign key[303] = 4557790;
assign key2[303] = 4878;
assign key3[303] = 0;
assign key[304] = 4548041;
assign key2[304] = 4870;
assign key3[304] = 0;
assign key[305] = 4538307;
assign key2[305] = 4863;
assign key3[305] = 0;
assign key[306] = 4528588;
assign key2[306] = 4856;
assign key3[306] = 0;
assign key[307] = 4518883;
assign key2[307] = 4848;
assign key3[307] = 0;
assign key[308] = 4509193;
assign key2[308] = 4841;
assign key3[308] = 0;
assign key[309] = 4499517;
assign key2[309] = 4834;
assign key3[309] = 0;
assign key[310] = 4489856;
assign key2[310] = 4827;
assign key3[310] = 0;
assign key[311] = 4480209;
assign key2[311] = 4819;
assign key3[311] = 0;
assign key[312] = 4470576;
assign key2[312] = 4812;
assign key3[312] = 0;
assign key[313] = 4460958;
assign key2[313] = 4805;
assign key3[313] = 0;
assign key[314] = 4451355;
assign key2[314] = 4798;
assign key3[314] = 0;
assign key[315] = 4441766;
assign key2[315] = 4791;
assign key3[315] = 0;
assign key[316] = 4432191;
assign key2[316] = 4783;
assign key3[316] = 0;
assign key[317] = 4422630;
assign key2[317] = 4776;
assign key3[317] = 0;
assign key[318] = 4413084;
assign key2[318] = 4769;
assign key3[318] = 0;
assign key[319] = 4403552;
assign key2[319] = 4762;
assign key3[319] = 0;
assign key[320] = 4394034;
assign key2[320] = 4755;
assign key3[320] = 0;
assign key[321] = 4384530;
assign key2[321] = 4748;
assign key3[321] = 0;
assign key[322] = 4375040;
assign key2[322] = 4741;
assign key3[322] = 0;
assign key[323] = 4365565;
assign key2[323] = 4734;
assign key3[323] = 0;
assign key[324] = 4356103;
assign key2[324] = 4727;
assign key3[324] = 0;
assign key[325] = 4346655;
assign key2[325] = 4720;
assign key3[325] = 0;
assign key[326] = 4337222;
assign key2[326] = 4713;
assign key3[326] = 0;
assign key[327] = 4327802;
assign key2[327] = 4706;
assign key3[327] = 0;
assign key[328] = 4318397;
assign key2[328] = 4699;
assign key3[328] = 0;
assign key[329] = 4309005;
assign key2[329] = 4692;
assign key3[329] = 0;
assign key[330] = 4299627;
assign key2[330] = 4685;
assign key3[330] = 0;
assign key[331] = 4290263;
assign key2[331] = 4678;
assign key3[331] = 0;
assign key[332] = 4280913;
assign key2[332] = 4671;
assign key3[332] = 0;
assign key[333] = 4271576;
assign key2[333] = 4664;
assign key3[333] = 0;
assign key[334] = 4262254;
assign key2[334] = 4657;
assign key3[334] = 0;
assign key[335] = 4252945;
assign key2[335] = 4651;
assign key3[335] = 0;
assign key[336] = 4243650;
assign key2[336] = 4644;
assign key3[336] = 0;
assign key[337] = 4234368;
assign key2[337] = 4637;
assign key3[337] = 0;
assign key[338] = 4225100;
assign key2[338] = 4630;
assign key3[338] = 0;
assign key[339] = 4215846;
assign key2[339] = 4623;
assign key3[339] = 0;
assign key[340] = 4206605;
assign key2[340] = 4617;
assign key3[340] = 0;
assign key[341] = 4197378;
assign key2[341] = 4610;
assign key3[341] = 0;
assign key[342] = 4188164;
assign key2[342] = 4603;
assign key3[342] = 0;
assign key[343] = 4178964;
assign key2[343] = 4596;
assign key3[343] = 0;
assign key[344] = 4169777;
assign key2[344] = 4590;
assign key3[344] = 0;
assign key[345] = 4160603;
assign key2[345] = 4583;
assign key3[345] = 0;
assign key[346] = 4151443;
assign key2[346] = 4576;
assign key3[346] = 0;
assign key[347] = 4142297;
assign key2[347] = 4569;
assign key3[347] = 0;
assign key[348] = 4133163;
assign key2[348] = 4563;
assign key3[348] = 0;
assign key[349] = 4124043;
assign key2[349] = 4556;
assign key3[349] = 0;
assign key[350] = 4114937;
assign key2[350] = 4550;
assign key3[350] = 0;
assign key[351] = 4105843;
assign key2[351] = 4543;
assign key3[351] = 0;
assign key[352] = 4096763;
assign key2[352] = 4536;
assign key3[352] = 0;
assign key[353] = 4087696;
assign key2[353] = 4530;
assign key3[353] = 0;
assign key[354] = 4078642;
assign key2[354] = 4523;
assign key3[354] = 0;
assign key[355] = 4069601;
assign key2[355] = 4517;
assign key3[355] = 0;
assign key[356] = 4060573;
assign key2[356] = 4510;
assign key3[356] = 0;
assign key[357] = 4051559;
assign key2[357] = 4504;
assign key3[357] = 0;
assign key[358] = 4042557;
assign key2[358] = 4497;
assign key3[358] = 0;
assign key[359] = 4033569;
assign key2[359] = 4491;
assign key3[359] = 0;
assign key[360] = 4024593;
assign key2[360] = 4484;
assign key3[360] = 0;
assign key[361] = 4015630;
assign key2[361] = 4478;
assign key3[361] = 0;
assign key[362] = 4006681;
assign key2[362] = 4471;
assign key3[362] = 0;
assign key[363] = 3997744;
assign key2[363] = 4465;
assign key3[363] = 0;
assign key[364] = 3988820;
assign key2[364] = 4458;
assign key3[364] = 0;
assign key[365] = 3979909;
assign key2[365] = 4452;
assign key3[365] = 0;
assign key[366] = 3971011;
assign key2[366] = 4445;
assign key3[366] = 0;
assign key[367] = 3962125;
assign key2[367] = 4439;
assign key3[367] = 0;
assign key[368] = 3953253;
assign key2[368] = 4433;
assign key3[368] = 0;
assign key[369] = 3944393;
assign key2[369] = 4426;
assign key3[369] = 0;
assign key[370] = 3935546;
assign key2[370] = 4420;
assign key3[370] = 0;
assign key[371] = 3926711;
assign key2[371] = 4414;
assign key3[371] = 0;
assign key[372] = 3917889;
assign key2[372] = 4407;
assign key3[372] = 0;
assign key[373] = 3909080;
assign key2[373] = 4401;
assign key3[373] = 0;
assign key[374] = 3900283;
assign key2[374] = 4395;
assign key3[374] = 0;
assign key[375] = 3891499;
assign key2[375] = 4388;
assign key3[375] = 0;
assign key[376] = 3882728;
assign key2[376] = 4382;
assign key3[376] = 0;
assign key[377] = 3873969;
assign key2[377] = 4376;
assign key3[377] = 0;
assign key[378] = 3865222;
assign key2[378] = 4370;
assign key3[378] = 0;
assign key[379] = 3856488;
assign key2[379] = 4363;
assign key3[379] = 0;
assign key[380] = 3847767;
assign key2[380] = 4357;
assign key3[380] = 0;
assign key[381] = 3839058;
assign key2[381] = 4351;
assign key3[381] = 0;
assign key[382] = 3830361;
assign key2[382] = 4345;
assign key3[382] = 0;
assign key[383] = 3821676;
assign key2[383] = 4339;
assign key3[383] = 0;
assign key[384] = 3813004;
assign key2[384] = 4332;
assign key3[384] = 0;
assign key[385] = 3804345;
assign key2[385] = 4326;
assign key3[385] = 0;
assign key[386] = 3795697;
assign key2[386] = 4320;
assign key3[386] = 0;
assign key[387] = 3787062;
assign key2[387] = 4314;
assign key3[387] = 0;
assign key[388] = 3778439;
assign key2[388] = 4308;
assign key3[388] = 0;
assign key[389] = 3769828;
assign key2[389] = 4302;
assign key3[389] = 0;
assign key[390] = 3761230;
assign key2[390] = 4296;
assign key3[390] = 0;
assign key[391] = 3752643;
assign key2[391] = 4290;
assign key3[391] = 0;
assign key[392] = 3744069;
assign key2[392] = 4284;
assign key3[392] = 0;
assign key[393] = 3735507;
assign key2[393] = 4278;
assign key3[393] = 0;
assign key[394] = 3726956;
assign key2[394] = 4272;
assign key3[394] = 0;
assign key[395] = 3718418;
assign key2[395] = 4266;
assign key3[395] = 0;
assign key[396] = 3709892;
assign key2[396] = 4260;
assign key3[396] = 0;
assign key[397] = 3701378;
assign key2[397] = 4254;
assign key3[397] = 0;
assign key[398] = 3692876;
assign key2[398] = 4248;
assign key3[398] = 0;
assign key[399] = 3684386;
assign key2[399] = 4242;
assign key3[399] = 0;
assign key[400] = 3675908;
assign key2[400] = 4236;
assign key3[400] = 0;
assign key[401] = 3667441;
assign key2[401] = 4230;
assign key3[401] = 0;
assign key[402] = 3658987;
assign key2[402] = 4224;
assign key3[402] = 0;
assign key[403] = 3650544;
assign key2[403] = 4218;
assign key3[403] = 0;
assign key[404] = 3642113;
assign key2[404] = 4212;
assign key3[404] = 0;
assign key[405] = 3633694;
assign key2[405] = 4206;
assign key3[405] = 0;
assign key[406] = 3625287;
assign key2[406] = 4200;
assign key3[406] = 0;
assign key[407] = 3616892;
assign key2[407] = 4194;
assign key3[407] = 0;
assign key[408] = 3608508;
assign key2[408] = 4188;
assign key3[408] = 0;
assign key[409] = 3600136;
assign key2[409] = 4183;
assign key3[409] = 0;
assign key[410] = 3591776;
assign key2[410] = 4177;
assign key3[410] = 0;
assign key[411] = 3583427;
assign key2[411] = 4171;
assign key3[411] = 0;
assign key[412] = 3575090;
assign key2[412] = 4165;
assign key3[412] = 0;
assign key[413] = 3566764;
assign key2[413] = 4159;
assign key3[413] = 0;
assign key[414] = 3558451;
assign key2[414] = 4154;
assign key3[414] = 0;
assign key[415] = 3550148;
assign key2[415] = 4148;
assign key3[415] = 0;
assign key[416] = 3541857;
assign key2[416] = 4142;
assign key3[416] = 0;
assign key[417] = 3533578;
assign key2[417] = 4136;
assign key3[417] = 0;
assign key[418] = 3525310;
assign key2[418] = 4131;
assign key3[418] = 0;
assign key[419] = 3517054;
assign key2[419] = 4125;
assign key3[419] = 0;
assign key[420] = 3508809;
assign key2[420] = 4119;
assign key3[420] = 0;
assign key[421] = 3500576;
assign key2[421] = 4113;
assign key3[421] = 0;
assign key[422] = 3492353;
assign key2[422] = 4108;
assign key3[422] = 0;
assign key[423] = 3484143;
assign key2[423] = 4102;
assign key3[423] = 0;
assign key[424] = 3475943;
assign key2[424] = 4096;
assign key3[424] = 0;
assign key[425] = 3467755;
assign key2[425] = 8182;
assign key3[425] = 1;
assign key[426] = 3459578;
assign key2[426] = 8171;
assign key3[426] = 1;
assign key[427] = 3451413;
assign key2[427] = 8159;
assign key3[427] = 1;
assign key[428] = 3443259;
assign key2[428] = 8148;
assign key3[428] = 1;
assign key[429] = 3435115;
assign key2[429] = 8137;
assign key3[429] = 1;
assign key[430] = 3426984;
assign key2[430] = 8126;
assign key3[430] = 1;
assign key[431] = 3418863;
assign key2[431] = 8115;
assign key3[431] = 1;
assign key[432] = 3410753;
assign key2[432] = 8103;
assign key3[432] = 1;
assign key[433] = 3402655;
assign key2[433] = 8092;
assign key3[433] = 1;
assign key[434] = 3394568;
assign key2[434] = 8081;
assign key3[434] = 1;
assign key[435] = 3386492;
assign key2[435] = 8070;
assign key3[435] = 1;
assign key[436] = 3378426;
assign key2[436] = 8059;
assign key3[436] = 1;
assign key[437] = 3370372;
assign key2[437] = 8048;
assign key3[437] = 1;
assign key[438] = 3362329;
assign key2[438] = 8037;
assign key3[438] = 1;
assign key[439] = 3354297;
assign key2[439] = 8026;
assign key3[439] = 1;
assign key[440] = 3346276;
assign key2[440] = 8015;
assign key3[440] = 1;
assign key[441] = 3338266;
assign key2[441] = 8004;
assign key3[441] = 1;
assign key[442] = 3330267;
assign key2[442] = 7993;
assign key3[442] = 1;
assign key[443] = 3322278;
assign key2[443] = 7982;
assign key3[443] = 1;
assign key[444] = 3314301;
assign key2[444] = 7972;
assign key3[444] = 1;
assign key[445] = 3306334;
assign key2[445] = 7961;
assign key3[445] = 1;
assign key[446] = 3298379;
assign key2[446] = 7950;
assign key3[446] = 1;
assign key[447] = 3290434;
assign key2[447] = 7939;
assign key3[447] = 1;
assign key[448] = 3282499;
assign key2[448] = 7928;
assign key3[448] = 1;
assign key[449] = 3274576;
assign key2[449] = 7917;
assign key3[449] = 1;
assign key[450] = 3266663;
assign key2[450] = 7907;
assign key3[450] = 1;
assign key[451] = 3258762;
assign key2[451] = 7896;
assign key3[451] = 1;
assign key[452] = 3250870;
assign key2[452] = 7885;
assign key3[452] = 1;
assign key[453] = 3242990;
assign key2[453] = 7875;
assign key3[453] = 1;
assign key[454] = 3235120;
assign key2[454] = 7864;
assign key3[454] = 1;
assign key[455] = 3227261;
assign key2[455] = 7853;
assign key3[455] = 1;
assign key[456] = 3219412;
assign key2[456] = 7843;
assign key3[456] = 1;
assign key[457] = 3211574;
assign key2[457] = 7832;
assign key3[457] = 1;
assign key[458] = 3203747;
assign key2[458] = 7822;
assign key3[458] = 1;
assign key[459] = 3195930;
assign key2[459] = 7811;
assign key3[459] = 1;
assign key[460] = 3188124;
assign key2[460] = 7801;
assign key3[460] = 1;
assign key[461] = 3180328;
assign key2[461] = 7790;
assign key3[461] = 1;
assign key[462] = 3172543;
assign key2[462] = 7780;
assign key3[462] = 1;
assign key[463] = 3164768;
assign key2[463] = 7769;
assign key3[463] = 1;
assign key[464] = 3157004;
assign key2[464] = 7759;
assign key3[464] = 1;
assign key[465] = 3149250;
assign key2[465] = 7748;
assign key3[465] = 1;
assign key[466] = 3141506;
assign key2[466] = 7738;
assign key3[466] = 1;
assign key[467] = 3133773;
assign key2[467] = 7727;
assign key3[467] = 1;
assign key[468] = 3126050;
assign key2[468] = 7717;
assign key3[468] = 1;
assign key[469] = 3118338;
assign key2[469] = 7707;
assign key3[469] = 1;
assign key[470] = 3110636;
assign key2[470] = 7696;
assign key3[470] = 1;
assign key[471] = 3102944;
assign key2[471] = 7686;
assign key3[471] = 1;
assign key[472] = 3095262;
assign key2[472] = 7676;
assign key3[472] = 1;
assign key[473] = 3087591;
assign key2[473] = 7666;
assign key3[473] = 1;
assign key[474] = 3079930;
assign key2[474] = 7655;
assign key3[474] = 1;
assign key[475] = 3072279;
assign key2[475] = 7645;
assign key3[475] = 1;
assign key[476] = 3064639;
assign key2[476] = 7635;
assign key3[476] = 1;
assign key[477] = 3057008;
assign key2[477] = 7625;
assign key3[477] = 1;
assign key[478] = 3049388;
assign key2[478] = 7615;
assign key3[478] = 1;
assign key[479] = 3041778;
assign key2[479] = 7605;
assign key3[479] = 1;
assign key[480] = 3034178;
assign key2[480] = 7594;
assign key3[480] = 1;
assign key[481] = 3026588;
assign key2[481] = 7584;
assign key3[481] = 1;
assign key[482] = 3019008;
assign key2[482] = 7574;
assign key3[482] = 1;
assign key[483] = 3011439;
assign key2[483] = 7564;
assign key3[483] = 1;
assign key[484] = 3003879;
assign key2[484] = 7554;
assign key3[484] = 1;
assign key[485] = 2996329;
assign key2[485] = 7544;
assign key3[485] = 1;
assign key[486] = 2988789;
assign key2[486] = 7534;
assign key3[486] = 1;
assign key[487] = 2981260;
assign key2[487] = 7524;
assign key3[487] = 1;
assign key[488] = 2973740;
assign key2[488] = 7514;
assign key3[488] = 1;
assign key[489] = 2966230;
assign key2[489] = 7504;
assign key3[489] = 1;
assign key[490] = 2958730;
assign key2[490] = 7494;
assign key3[490] = 1;
assign key[491] = 2951240;
assign key2[491] = 7485;
assign key3[491] = 1;
assign key[492] = 2943760;
assign key2[492] = 7475;
assign key3[492] = 1;
assign key[493] = 2936290;
assign key2[493] = 7465;
assign key3[493] = 1;
assign key[494] = 2928829;
assign key2[494] = 7455;
assign key3[494] = 1;
assign key[495] = 2921379;
assign key2[495] = 7445;
assign key3[495] = 1;
assign key[496] = 2913938;
assign key2[496] = 7435;
assign key3[496] = 1;
assign key[497] = 2906507;
assign key2[497] = 7426;
assign key3[497] = 1;
assign key[498] = 2899086;
assign key2[498] = 7416;
assign key3[498] = 1;
assign key[499] = 2891674;
assign key2[499] = 7406;
assign key3[499] = 1;
assign key[500] = 2884273;
assign key2[500] = 7396;
assign key3[500] = 1;
assign key[501] = 2876881;
assign key2[501] = 7387;
assign key3[501] = 1;
assign key[502] = 2869498;
assign key2[502] = 7377;
assign key3[502] = 1;
assign key[503] = 2862126;
assign key2[503] = 7367;
assign key3[503] = 1;
assign key[504] = 2854762;
assign key2[504] = 7358;
assign key3[504] = 1;
assign key[505] = 2847409;
assign key2[505] = 7348;
assign key3[505] = 1;
assign key[506] = 2840065;
assign key2[506] = 7339;
assign key3[506] = 1;
assign key[507] = 2832731;
assign key2[507] = 7329;
assign key3[507] = 1;
assign key[508] = 2825406;
assign key2[508] = 7319;
assign key3[508] = 1;
assign key[509] = 2818091;
assign key2[509] = 7310;
assign key3[509] = 1;
assign key[510] = 2810786;
assign key2[510] = 7300;
assign key3[510] = 1;
assign key[511] = 2803490;
assign key2[511] = 7291;
assign key3[511] = 1;
assign key[512] = 2796203;
assign key2[512] = 7281;
assign key3[512] = 1;
assign key[513] = 2788926;
assign key2[513] = 7272;
assign key3[513] = 1;
assign key[514] = 2781659;
assign key2[514] = 7262;
assign key3[514] = 1;
assign key[515] = 2774401;
assign key2[515] = 7253;
assign key3[515] = 1;
assign key[516] = 2767152;
assign key2[516] = 7243;
assign key3[516] = 1;
assign key[517] = 2759912;
assign key2[517] = 7234;
assign key3[517] = 1;
assign key[518] = 2752683;
assign key2[518] = 7225;
assign key3[518] = 1;
assign key[519] = 2745462;
assign key2[519] = 7215;
assign key3[519] = 1;
assign key[520] = 2738251;
assign key2[520] = 7206;
assign key3[520] = 1;
assign key[521] = 2731049;
assign key2[521] = 7197;
assign key3[521] = 1;
assign key[522] = 2723856;
assign key2[522] = 7187;
assign key3[522] = 1;
assign key[523] = 2716673;
assign key2[523] = 7178;
assign key3[523] = 1;
assign key[524] = 2709499;
assign key2[524] = 7169;
assign key3[524] = 1;
assign key[525] = 2702335;
assign key2[525] = 7160;
assign key3[525] = 1;
assign key[526] = 2695179;
assign key2[526] = 7150;
assign key3[526] = 1;
assign key[527] = 2688033;
assign key2[527] = 7141;
assign key3[527] = 1;
assign key[528] = 2680896;
assign key2[528] = 7132;
assign key3[528] = 1;
assign key[529] = 2673768;
assign key2[529] = 7123;
assign key3[529] = 1;
assign key[530] = 2666649;
assign key2[530] = 7114;
assign key3[530] = 1;
assign key[531] = 2659540;
assign key2[531] = 7104;
assign key3[531] = 1;
assign key[532] = 2652440;
assign key2[532] = 7095;
assign key3[532] = 1;
assign key[533] = 2645348;
assign key2[533] = 7086;
assign key3[533] = 1;
assign key[534] = 2638266;
assign key2[534] = 7077;
assign key3[534] = 1;
assign key[535] = 2631193;
assign key2[535] = 7068;
assign key3[535] = 1;
assign key[536] = 2624129;
assign key2[536] = 7059;
assign key3[536] = 1;
assign key[537] = 2617074;
assign key2[537] = 7050;
assign key3[537] = 1;
assign key[538] = 2610028;
assign key2[538] = 7041;
assign key3[538] = 1;
assign key[539] = 2602992;
assign key2[539] = 7032;
assign key3[539] = 1;
assign key[540] = 2595964;
assign key2[540] = 7023;
assign key3[540] = 1;
assign key[541] = 2588945;
assign key2[541] = 7014;
assign key3[541] = 1;
assign key[542] = 2581935;
assign key2[542] = 7005;
assign key3[542] = 1;
assign key[543] = 2574934;
assign key2[543] = 6996;
assign key3[543] = 1;
assign key[544] = 2567942;
assign key2[544] = 6987;
assign key3[544] = 1;
assign key[545] = 2560959;
assign key2[545] = 6978;
assign key3[545] = 1;
assign key[546] = 2553984;
assign key2[546] = 6969;
assign key3[546] = 1;
assign key[547] = 2547019;
assign key2[547] = 6960;
assign key3[547] = 1;
assign key[548] = 2540063;
assign key2[548] = 6952;
assign key3[548] = 1;
assign key[549] = 2533115;
assign key2[549] = 6943;
assign key3[549] = 1;
assign key[550] = 2526176;
assign key2[550] = 6934;
assign key3[550] = 1;
assign key[551] = 2519246;
assign key2[551] = 6925;
assign key3[551] = 1;
assign key[552] = 2512325;
assign key2[552] = 6916;
assign key3[552] = 1;
assign key[553] = 2505412;
assign key2[553] = 6908;
assign key3[553] = 1;
assign key[554] = 2498509;
assign key2[554] = 6899;
assign key3[554] = 1;
assign key[555] = 2491614;
assign key2[555] = 6890;
assign key3[555] = 1;
assign key[556] = 2484727;
assign key2[556] = 6881;
assign key3[556] = 1;
assign key[557] = 2477850;
assign key2[557] = 6873;
assign key3[557] = 1;
assign key[558] = 2470981;
assign key2[558] = 6864;
assign key3[558] = 1;
assign key[559] = 2464121;
assign key2[559] = 6855;
assign key3[559] = 1;
assign key[560] = 2457270;
assign key2[560] = 6847;
assign key3[560] = 1;
assign key[561] = 2450427;
assign key2[561] = 6838;
assign key3[561] = 1;
assign key[562] = 2443593;
assign key2[562] = 6829;
assign key3[562] = 1;
assign key[563] = 2436767;
assign key2[563] = 6821;
assign key3[563] = 1;
assign key[564] = 2429950;
assign key2[564] = 6812;
assign key3[564] = 1;
assign key[565] = 2423142;
assign key2[565] = 6804;
assign key3[565] = 1;
assign key[566] = 2416342;
assign key2[566] = 6795;
assign key3[566] = 1;
assign key[567] = 2409550;
assign key2[567] = 6787;
assign key3[567] = 1;
assign key[568] = 2402768;
assign key2[568] = 6778;
assign key3[568] = 1;
assign key[569] = 2395993;
assign key2[569] = 6769;
assign key3[569] = 1;
assign key[570] = 2389228;
assign key2[570] = 6761;
assign key3[570] = 1;
assign key[571] = 2382470;
assign key2[571] = 6753;
assign key3[571] = 1;
assign key[572] = 2375722;
assign key2[572] = 6744;
assign key3[572] = 1;
assign key[573] = 2368981;
assign key2[573] = 6736;
assign key3[573] = 1;
assign key[574] = 2362249;
assign key2[574] = 6727;
assign key3[574] = 1;
assign key[575] = 2355526;
assign key2[575] = 6719;
assign key3[575] = 1;
assign key[576] = 2348811;
assign key2[576] = 6710;
assign key3[576] = 1;
assign key[577] = 2342104;
assign key2[577] = 6702;
assign key3[577] = 1;
assign key[578] = 2335406;
assign key2[578] = 6694;
assign key3[578] = 1;
assign key[579] = 2328716;
assign key2[579] = 6685;
assign key3[579] = 1;
assign key[580] = 2322034;
assign key2[580] = 6677;
assign key3[580] = 1;
assign key[581] = 2315361;
assign key2[581] = 6669;
assign key3[581] = 1;
assign key[582] = 2308696;
assign key2[582] = 6660;
assign key3[582] = 1;
assign key[583] = 2302039;
assign key2[583] = 6652;
assign key3[583] = 1;
assign key[584] = 2295391;
assign key2[584] = 6644;
assign key3[584] = 1;
assign key[585] = 2288751;
assign key2[585] = 6636;
assign key3[585] = 1;
assign key[586] = 2282119;
assign key2[586] = 6627;
assign key3[586] = 1;
assign key[587] = 2275495;
assign key2[587] = 6619;
assign key3[587] = 1;
assign key[588] = 2268880;
assign key2[588] = 6611;
assign key3[588] = 1;
assign key[589] = 2262272;
assign key2[589] = 6603;
assign key3[589] = 1;
assign key[590] = 2255673;
assign key2[590] = 6594;
assign key3[590] = 1;
assign key[591] = 2249082;
assign key2[591] = 6586;
assign key3[591] = 1;
assign key[592] = 2242500;
assign key2[592] = 6578;
assign key3[592] = 1;
assign key[593] = 2235925;
assign key2[593] = 6570;
assign key3[593] = 1;
assign key[594] = 2229359;
assign key2[594] = 6562;
assign key3[594] = 1;
assign key[595] = 2222800;
assign key2[595] = 6554;
assign key3[595] = 1;
assign key[596] = 2216250;
assign key2[596] = 6546;
assign key3[596] = 1;
assign key[597] = 2209708;
assign key2[597] = 6538;
assign key3[597] = 1;
assign key[598] = 2203174;
assign key2[598] = 6530;
assign key3[598] = 1;
assign key[599] = 2196648;
assign key2[599] = 6522;
assign key3[599] = 1;
assign key[600] = 2190130;
assign key2[600] = 6514;
assign key3[600] = 1;
assign key[601] = 2183620;
assign key2[601] = 6505;
assign key3[601] = 1;
assign key[602] = 2177118;
assign key2[602] = 6497;
assign key3[602] = 1;
assign key[603] = 2170624;
assign key2[603] = 6490;
assign key3[603] = 1;
assign key[604] = 2164138;
assign key2[604] = 6482;
assign key3[604] = 1;
assign key[605] = 2157660;
assign key2[605] = 6474;
assign key3[605] = 1;
assign key[606] = 2151190;
assign key2[606] = 6466;
assign key3[606] = 1;
assign key[607] = 2144727;
assign key2[607] = 6458;
assign key3[607] = 1;
assign key[608] = 2138273;
assign key2[608] = 6450;
assign key3[608] = 1;
assign key[609] = 2131827;
assign key2[609] = 6442;
assign key3[609] = 1;
assign key[610] = 2125388;
assign key2[610] = 6434;
assign key3[610] = 1;
assign key[611] = 2118958;
assign key2[611] = 6426;
assign key3[611] = 1;
assign key[612] = 2112535;
assign key2[612] = 6418;
assign key3[612] = 1;
assign key[613] = 2106120;
assign key2[613] = 6410;
assign key3[613] = 1;
assign key[614] = 2099713;
assign key2[614] = 6403;
assign key3[614] = 1;
assign key[615] = 2093314;
assign key2[615] = 6395;
assign key3[615] = 1;
assign key[616] = 2086922;
assign key2[616] = 6387;
assign key3[616] = 1;
assign key[617] = 2080539;
assign key2[617] = 6379;
assign key3[617] = 1;
assign key[618] = 2074163;
assign key2[618] = 6371;
assign key3[618] = 1;
assign key[619] = 2067795;
assign key2[619] = 6364;
assign key3[619] = 1;
assign key[620] = 2061435;
assign key2[620] = 6356;
assign key3[620] = 1;
assign key[621] = 2055082;
assign key2[621] = 6348;
assign key3[621] = 1;
assign key[622] = 2048737;
assign key2[622] = 6341;
assign key3[622] = 1;
assign key[623] = 2042400;
assign key2[623] = 6333;
assign key3[623] = 1;
assign key[624] = 2036070;
assign key2[624] = 6325;
assign key3[624] = 1;
assign key[625] = 2029749;
assign key2[625] = 6317;
assign key3[625] = 1;
assign key[626] = 2023434;
assign key2[626] = 6310;
assign key3[626] = 1;
assign key[627] = 2017128;
assign key2[627] = 6302;
assign key3[627] = 1;
assign key[628] = 2010829;
assign key2[628] = 6295;
assign key3[628] = 1;
assign key[629] = 2004538;
assign key2[629] = 6287;
assign key3[629] = 1;
assign key[630] = 1998254;
assign key2[630] = 6279;
assign key3[630] = 1;
assign key[631] = 1991978;
assign key2[631] = 6272;
assign key3[631] = 1;
assign key[632] = 1985710;
assign key2[632] = 6264;
assign key3[632] = 1;
assign key[633] = 1979449;
assign key2[633] = 6257;
assign key3[633] = 1;
assign key[634] = 1973195;
assign key2[634] = 6249;
assign key3[634] = 1;
assign key[635] = 1966950;
assign key2[635] = 6242;
assign key3[635] = 1;
assign key[636] = 1960711;
assign key2[636] = 6234;
assign key3[636] = 1;
assign key[637] = 1954480;
assign key2[637] = 6227;
assign key3[637] = 1;
assign key[638] = 1948257;
assign key2[638] = 6219;
assign key3[638] = 1;
assign key[639] = 1942041;
assign key2[639] = 6212;
assign key3[639] = 1;
assign key[640] = 1935833;
assign key2[640] = 6204;
assign key3[640] = 1;
assign key[641] = 1929632;
assign key2[641] = 6197;
assign key3[641] = 1;
assign key[642] = 1923439;
assign key2[642] = 6189;
assign key3[642] = 1;
assign key[643] = 1917253;
assign key2[643] = 6182;
assign key3[643] = 1;
assign key[644] = 1911074;
assign key2[644] = 6174;
assign key3[644] = 1;
assign key[645] = 1904903;
assign key2[645] = 6167;
assign key3[645] = 1;
assign key[646] = 1898739;
assign key2[646] = 6160;
assign key3[646] = 1;
assign key[647] = 1892583;
assign key2[647] = 6152;
assign key3[647] = 1;
assign key[648] = 1886434;
assign key2[648] = 6145;
assign key3[648] = 1;
assign key[649] = 1880292;
assign key2[649] = 6138;
assign key3[649] = 1;
assign key[650] = 1874158;
assign key2[650] = 6130;
assign key3[650] = 1;
assign key[651] = 1868031;
assign key2[651] = 6123;
assign key3[651] = 1;
assign key[652] = 1861911;
assign key2[652] = 6116;
assign key3[652] = 1;
assign key[653] = 1855799;
assign key2[653] = 6108;
assign key3[653] = 1;
assign key[654] = 1849694;
assign key2[654] = 6101;
assign key3[654] = 1;
assign key[655] = 1843596;
assign key2[655] = 6094;
assign key3[655] = 1;
assign key[656] = 1837505;
assign key2[656] = 6086;
assign key3[656] = 1;
assign key[657] = 1831422;
assign key2[657] = 6079;
assign key3[657] = 1;
assign key[658] = 1825346;
assign key2[658] = 6072;
assign key3[658] = 1;
assign key[659] = 1819277;
assign key2[659] = 6065;
assign key3[659] = 1;
assign key[660] = 1813215;
assign key2[660] = 6058;
assign key3[660] = 1;
assign key[661] = 1807161;
assign key2[661] = 6050;
assign key3[661] = 1;
assign key[662] = 1801113;
assign key2[662] = 6043;
assign key3[662] = 1;
assign key[663] = 1795073;
assign key2[663] = 6036;
assign key3[663] = 1;
assign key[664] = 1789040;
assign key2[664] = 6029;
assign key3[664] = 1;
assign key[665] = 1783014;
assign key2[665] = 6022;
assign key3[665] = 1;
assign key[666] = 1776996;
assign key2[666] = 6015;
assign key3[666] = 1;
assign key[667] = 1770984;
assign key2[667] = 6008;
assign key3[667] = 1;
assign key[668] = 1764979;
assign key2[668] = 6000;
assign key3[668] = 1;
assign key[669] = 1758982;
assign key2[669] = 5993;
assign key3[669] = 1;
assign key[670] = 1752992;
assign key2[670] = 5986;
assign key3[670] = 1;
assign key[671] = 1747008;
assign key2[671] = 5979;
assign key3[671] = 1;
assign key[672] = 1741032;
assign key2[672] = 5972;
assign key3[672] = 1;
assign key[673] = 1735063;
assign key2[673] = 5965;
assign key3[673] = 1;
assign key[674] = 1729101;
assign key2[674] = 5958;
assign key3[674] = 1;
assign key[675] = 1723146;
assign key2[675] = 5951;
assign key3[675] = 1;
assign key[676] = 1717198;
assign key2[676] = 5944;
assign key3[676] = 1;
assign key[677] = 1711257;
assign key2[677] = 5937;
assign key3[677] = 1;
assign key[678] = 1705323;
assign key2[678] = 5930;
assign key3[678] = 1;
assign key[679] = 1699395;
assign key2[679] = 5923;
assign key3[679] = 1;
assign key[680] = 1693475;
assign key2[680] = 5916;
assign key3[680] = 1;
assign key[681] = 1687562;
assign key2[681] = 5909;
assign key3[681] = 1;
assign key[682] = 1681656;
assign key2[682] = 5902;
assign key3[682] = 1;
assign key[683] = 1675756;
assign key2[683] = 5895;
assign key3[683] = 1;
assign key[684] = 1669864;
assign key2[684] = 5889;
assign key3[684] = 1;
assign key[685] = 1663978;
assign key2[685] = 5882;
assign key3[685] = 1;
assign key[686] = 1658100;
assign key2[686] = 5875;
assign key3[686] = 1;
assign key[687] = 1652228;
assign key2[687] = 5868;
assign key3[687] = 1;
assign key[688] = 1646363;
assign key2[688] = 5861;
assign key3[688] = 1;
assign key[689] = 1640505;
assign key2[689] = 5854;
assign key3[689] = 1;
assign key[690] = 1634653;
assign key2[690] = 5847;
assign key3[690] = 1;
assign key[691] = 1628809;
assign key2[691] = 5841;
assign key3[691] = 1;
assign key[692] = 1622971;
assign key2[692] = 5834;
assign key3[692] = 1;
assign key[693] = 1617140;
assign key2[693] = 5827;
assign key3[693] = 1;
assign key[694] = 1611316;
assign key2[694] = 5820;
assign key3[694] = 1;
assign key[695] = 1605499;
assign key2[695] = 5813;
assign key3[695] = 1;
assign key[696] = 1599688;
assign key2[696] = 5807;
assign key3[696] = 1;
assign key[697] = 1593885;
assign key2[697] = 5800;
assign key3[697] = 1;
assign key[698] = 1588088;
assign key2[698] = 5793;
assign key3[698] = 1;
assign key[699] = 1582297;
assign key2[699] = 5786;
assign key3[699] = 1;
assign key[700] = 1576514;
assign key2[700] = 5780;
assign key3[700] = 1;
assign key[701] = 1570737;
assign key2[701] = 5773;
assign key3[701] = 1;
assign key[702] = 1564967;
assign key2[702] = 5766;
assign key3[702] = 1;
assign key[703] = 1559203;
assign key2[703] = 5760;
assign key3[703] = 1;
assign key[704] = 1553446;
assign key2[704] = 5753;
assign key3[704] = 1;
assign key[705] = 1547696;
assign key2[705] = 5746;
assign key3[705] = 1;
assign key[706] = 1541953;
assign key2[706] = 5740;
assign key3[706] = 1;
assign key[707] = 1536216;
assign key2[707] = 5733;
assign key3[707] = 1;
assign key[708] = 1530485;
assign key2[708] = 5726;
assign key3[708] = 1;
assign key[709] = 1524762;
assign key2[709] = 5720;
assign key3[709] = 1;
assign key[710] = 1519045;
assign key2[710] = 5713;
assign key3[710] = 1;
assign key[711] = 1513334;
assign key2[711] = 5707;
assign key3[711] = 1;
assign key[712] = 1507630;
assign key2[712] = 5700;
assign key3[712] = 1;
assign key[713] = 1501933;
assign key2[713] = 5694;
assign key3[713] = 1;
assign key[714] = 1496242;
assign key2[714] = 5687;
assign key3[714] = 1;
assign key[715] = 1490558;
assign key2[715] = 5680;
assign key3[715] = 1;
assign key[716] = 1484880;
assign key2[716] = 5674;
assign key3[716] = 1;
assign key[717] = 1479209;
assign key2[717] = 5667;
assign key3[717] = 1;
assign key[718] = 1473545;
assign key2[718] = 5661;
assign key3[718] = 1;
assign key[719] = 1467886;
assign key2[719] = 5654;
assign key3[719] = 1;
assign key[720] = 1462235;
assign key2[720] = 5648;
assign key3[720] = 1;
assign key[721] = 1456590;
assign key2[721] = 5641;
assign key3[721] = 1;
assign key[722] = 1450951;
assign key2[722] = 5635;
assign key3[722] = 1;
assign key[723] = 1445319;
assign key2[723] = 5629;
assign key3[723] = 1;
assign key[724] = 1439693;
assign key2[724] = 5622;
assign key3[724] = 1;
assign key[725] = 1434073;
assign key2[725] = 5616;
assign key3[725] = 1;
assign key[726] = 1428461;
assign key2[726] = 5609;
assign key3[726] = 1;
assign key[727] = 1422854;
assign key2[727] = 5603;
assign key3[727] = 1;
assign key[728] = 1417254;
assign key2[728] = 5596;
assign key3[728] = 1;
assign key[729] = 1411660;
assign key2[729] = 5590;
assign key3[729] = 1;
assign key[730] = 1406073;
assign key2[730] = 5584;
assign key3[730] = 1;
assign key[731] = 1400492;
assign key2[731] = 5577;
assign key3[731] = 1;
assign key[732] = 1394917;
assign key2[732] = 5571;
assign key3[732] = 1;
assign key[733] = 1389349;
assign key2[733] = 5565;
assign key3[733] = 1;
assign key[734] = 1383787;
assign key2[734] = 5558;
assign key3[734] = 1;
assign key[735] = 1378231;
assign key2[735] = 5552;
assign key3[735] = 1;
assign key[736] = 1372682;
assign key2[736] = 5546;
assign key3[736] = 1;
assign key[737] = 1367139;
assign key2[737] = 5539;
assign key3[737] = 1;
assign key[738] = 1361602;
assign key2[738] = 5533;
assign key3[738] = 1;
assign key[739] = 1356071;
assign key2[739] = 5527;
assign key3[739] = 1;
assign key[740] = 1350547;
assign key2[740] = 5521;
assign key3[740] = 1;
assign key[741] = 1345029;
assign key2[741] = 5514;
assign key3[741] = 1;
assign key[742] = 1339518;
assign key2[742] = 5508;
assign key3[742] = 1;
assign key[743] = 1334012;
assign key2[743] = 5502;
assign key3[743] = 1;
assign key[744] = 1328513;
assign key2[744] = 5496;
assign key3[744] = 1;
assign key[745] = 1323020;
assign key2[745] = 5489;
assign key3[745] = 1;
assign key[746] = 1317533;
assign key2[746] = 5483;
assign key3[746] = 1;
assign key[747] = 1312053;
assign key2[747] = 5477;
assign key3[747] = 1;
assign key[748] = 1306578;
assign key2[748] = 5471;
assign key3[748] = 1;
assign key[749] = 1301110;
assign key2[749] = 5465;
assign key3[749] = 1;
assign key[750] = 1295648;
assign key2[750] = 5458;
assign key3[750] = 1;
assign key[751] = 1290192;
assign key2[751] = 5452;
assign key3[751] = 1;
assign key[752] = 1284742;
assign key2[752] = 5446;
assign key3[752] = 1;
assign key[753] = 1279299;
assign key2[753] = 5440;
assign key3[753] = 1;
assign key[754] = 1273861;
assign key2[754] = 5434;
assign key3[754] = 1;
assign key[755] = 1268430;
assign key2[755] = 5428;
assign key3[755] = 1;
assign key[756] = 1263004;
assign key2[756] = 5422;
assign key3[756] = 1;
assign key[757] = 1257585;
assign key2[757] = 5416;
assign key3[757] = 1;
assign key[758] = 1252172;
assign key2[758] = 5410;
assign key3[758] = 1;
assign key[759] = 1246765;
assign key2[759] = 5404;
assign key3[759] = 1;
assign key[760] = 1241364;
assign key2[760] = 5397;
assign key3[760] = 1;
assign key[761] = 1235969;
assign key2[761] = 5391;
assign key3[761] = 1;
assign key[762] = 1230580;
assign key2[762] = 5385;
assign key3[762] = 1;
assign key[763] = 1225197;
assign key2[763] = 5379;
assign key3[763] = 1;
assign key[764] = 1219820;
assign key2[764] = 5373;
assign key3[764] = 1;
assign key[765] = 1214449;
assign key2[765] = 5367;
assign key3[765] = 1;
assign key[766] = 1209085;
assign key2[766] = 5361;
assign key3[766] = 1;
assign key[767] = 1203726;
assign key2[767] = 5355;
assign key3[767] = 1;
assign key[768] = 1198373;
assign key2[768] = 5349;
assign key3[768] = 1;
assign key[769] = 1193026;
assign key2[769] = 5343;
assign key3[769] = 1;
assign key[770] = 1187685;
assign key2[770] = 5337;
assign key3[770] = 1;
assign key[771] = 1182350;
assign key2[771] = 5332;
assign key3[771] = 1;
assign key[772] = 1177021;
assign key2[772] = 5326;
assign key3[772] = 1;
assign key[773] = 1171698;
assign key2[773] = 5320;
assign key3[773] = 1;
assign key[774] = 1166381;
assign key2[774] = 5314;
assign key3[774] = 1;
assign key[775] = 1161070;
assign key2[775] = 5308;
assign key3[775] = 1;
assign key[776] = 1155764;
assign key2[776] = 5302;
assign key3[776] = 1;
assign key[777] = 1150465;
assign key2[777] = 5296;
assign key3[777] = 1;
assign key[778] = 1145171;
assign key2[778] = 5290;
assign key3[778] = 1;
assign key[779] = 1139883;
assign key2[779] = 5284;
assign key3[779] = 1;
assign key[780] = 1134601;
assign key2[780] = 5278;
assign key3[780] = 1;
assign key[781] = 1129325;
assign key2[781] = 5273;
assign key3[781] = 1;
assign key[782] = 1124055;
assign key2[782] = 5267;
assign key3[782] = 1;
assign key[783] = 1118791;
assign key2[783] = 5261;
assign key3[783] = 1;
assign key[784] = 1113532;
assign key2[784] = 5255;
assign key3[784] = 1;
assign key[785] = 1108280;
assign key2[785] = 5249;
assign key3[785] = 1;
assign key[786] = 1103033;
assign key2[786] = 5244;
assign key3[786] = 1;
assign key[787] = 1097792;
assign key2[787] = 5238;
assign key3[787] = 1;
assign key[788] = 1092556;
assign key2[788] = 5232;
assign key3[788] = 1;
assign key[789] = 1087327;
assign key2[789] = 5226;
assign key3[789] = 1;
assign key[790] = 1082103;
assign key2[790] = 5220;
assign key3[790] = 1;
assign key[791] = 1076885;
assign key2[791] = 5215;
assign key3[791] = 1;
assign key[792] = 1071673;
assign key2[792] = 5209;
assign key3[792] = 1;
assign key[793] = 1066466;
assign key2[793] = 5203;
assign key3[793] = 1;
assign key[794] = 1061265;
assign key2[794] = 5197;
assign key3[794] = 1;
assign key[795] = 1056070;
assign key2[795] = 5192;
assign key3[795] = 1;
assign key[796] = 1050881;
assign key2[796] = 5186;
assign key3[796] = 1;
assign key[797] = 1045697;
assign key2[797] = 5180;
assign key3[797] = 1;
assign key[798] = 1040519;
assign key2[798] = 5175;
assign key3[798] = 1;
assign key[799] = 1035347;
assign key2[799] = 5169;
assign key3[799] = 1;
assign key[800] = 1030180;
assign key2[800] = 5163;
assign key3[800] = 1;
assign key[801] = 1025019;
assign key2[801] = 5158;
assign key3[801] = 1;
assign key[802] = 1019864;
assign key2[802] = 5152;
assign key3[802] = 1;
assign key[803] = 1014714;
assign key2[803] = 5146;
assign key3[803] = 1;
assign key[804] = 1009570;
assign key2[804] = 5141;
assign key3[804] = 1;
assign key[805] = 1004432;
assign key2[805] = 5135;
assign key3[805] = 1;
assign key[806] = 999299;
assign key2[806] = 5130;
assign key3[806] = 1;
assign key[807] = 994172;
assign key2[807] = 5124;
assign key3[807] = 1;
assign key[808] = 989050;
assign key2[808] = 5118;
assign key3[808] = 1;
assign key[809] = 983934;
assign key2[809] = 5113;
assign key3[809] = 1;
assign key[810] = 978824;
assign key2[810] = 5107;
assign key3[810] = 1;
assign key[811] = 973719;
assign key2[811] = 5102;
assign key3[811] = 1;
assign key[812] = 968620;
assign key2[812] = 5096;
assign key3[812] = 1;
assign key[813] = 963526;
assign key2[813] = 5090;
assign key3[813] = 1;
assign key[814] = 958438;
assign key2[814] = 5085;
assign key3[814] = 1;
assign key[815] = 953355;
assign key2[815] = 5079;
assign key3[815] = 1;
assign key[816] = 948278;
assign key2[816] = 5074;
assign key3[816] = 1;
assign key[817] = 943206;
assign key2[817] = 5068;
assign key3[817] = 1;
assign key[818] = 938140;
assign key2[818] = 5063;
assign key3[818] = 1;
assign key[819] = 933079;
assign key2[819] = 5057;
assign key3[819] = 1;
assign key[820] = 928024;
assign key2[820] = 5052;
assign key3[820] = 1;
assign key[821] = 922975;
assign key2[821] = 5046;
assign key3[821] = 1;
assign key[822] = 917930;
assign key2[822] = 5041;
assign key3[822] = 1;
assign key[823] = 912892;
assign key2[823] = 5036;
assign key3[823] = 1;
assign key[824] = 907858;
assign key2[824] = 5030;
assign key3[824] = 1;
assign key[825] = 902831;
assign key2[825] = 5025;
assign key3[825] = 1;
assign key[826] = 897808;
assign key2[826] = 5019;
assign key3[826] = 1;
assign key[827] = 892791;
assign key2[827] = 5014;
assign key3[827] = 1;
assign key[828] = 887780;
assign key2[828] = 5008;
assign key3[828] = 1;
assign key[829] = 882773;
assign key2[829] = 5003;
assign key3[829] = 1;
assign key[830] = 877773;
assign key2[830] = 4998;
assign key3[830] = 1;
assign key[831] = 872777;
assign key2[831] = 4992;
assign key3[831] = 1;
assign key[832] = 867787;
assign key2[832] = 4987;
assign key3[832] = 1;
assign key[833] = 862803;
assign key2[833] = 4981;
assign key3[833] = 1;
assign key[834] = 857824;
assign key2[834] = 4976;
assign key3[834] = 1;
assign key[835] = 852850;
assign key2[835] = 4971;
assign key3[835] = 1;
assign key[836] = 847881;
assign key2[836] = 4965;
assign key3[836] = 1;
assign key[837] = 842918;
assign key2[837] = 4960;
assign key3[837] = 1;
assign key[838] = 837960;
assign key2[838] = 4955;
assign key3[838] = 1;
assign key[839] = 833008;
assign key2[839] = 4949;
assign key3[839] = 1;
assign key[840] = 828060;
assign key2[840] = 4944;
assign key3[840] = 1;
assign key[841] = 823118;
assign key2[841] = 4939;
assign key3[841] = 1;
assign key[842] = 818182;
assign key2[842] = 4933;
assign key3[842] = 1;
assign key[843] = 813250;
assign key2[843] = 4928;
assign key3[843] = 1;
assign key[844] = 808324;
assign key2[844] = 4923;
assign key3[844] = 1;
assign key[845] = 803404;
assign key2[845] = 4918;
assign key3[845] = 1;
assign key[846] = 798488;
assign key2[846] = 4912;
assign key3[846] = 1;
assign key[847] = 793578;
assign key2[847] = 4907;
assign key3[847] = 1;
assign key[848] = 788673;
assign key2[848] = 4902;
assign key3[848] = 1;
assign key[849] = 783773;
assign key2[849] = 4897;
assign key3[849] = 1;
assign key[850] = 778879;
assign key2[850] = 4891;
assign key3[850] = 1;
assign key[851] = 773989;
assign key2[851] = 4886;
assign key3[851] = 1;
assign key[852] = 769105;
assign key2[852] = 4881;
assign key3[852] = 1;
assign key[853] = 764226;
assign key2[853] = 4876;
assign key3[853] = 1;
assign key[854] = 759352;
assign key2[854] = 4871;
assign key3[854] = 1;
assign key[855] = 754484;
assign key2[855] = 4865;
assign key3[855] = 1;
assign key[856] = 749621;
assign key2[856] = 4860;
assign key3[856] = 1;
assign key[857] = 744762;
assign key2[857] = 4855;
assign key3[857] = 1;
assign key[858] = 739909;
assign key2[858] = 4850;
assign key3[858] = 1;
assign key[859] = 735062;
assign key2[859] = 4845;
assign key3[859] = 1;
assign key[860] = 730219;
assign key2[860] = 4840;
assign key3[860] = 1;
assign key[861] = 725381;
assign key2[861] = 4835;
assign key3[861] = 1;
assign key[862] = 720549;
assign key2[862] = 4829;
assign key3[862] = 1;
assign key[863] = 715722;
assign key2[863] = 4824;
assign key3[863] = 1;
assign key[864] = 710899;
assign key2[864] = 4819;
assign key3[864] = 1;
assign key[865] = 706082;
assign key2[865] = 4814;
assign key3[865] = 1;
assign key[866] = 701270;
assign key2[866] = 4809;
assign key3[866] = 1;
assign key[867] = 696463;
assign key2[867] = 4804;
assign key3[867] = 1;
assign key[868] = 691661;
assign key2[868] = 4799;
assign key3[868] = 1;
assign key[869] = 686865;
assign key2[869] = 4794;
assign key3[869] = 1;
assign key[870] = 682073;
assign key2[870] = 4789;
assign key3[870] = 1;
assign key[871] = 677286;
assign key2[871] = 4784;
assign key3[871] = 1;
assign key[872] = 672505;
assign key2[872] = 4779;
assign key3[872] = 1;
assign key[873] = 667728;
assign key2[873] = 4774;
assign key3[873] = 1;
assign key[874] = 662957;
assign key2[874] = 4769;
assign key3[874] = 1;
assign key[875] = 658190;
assign key2[875] = 4763;
assign key3[875] = 1;
assign key[876] = 653429;
assign key2[876] = 4758;
assign key3[876] = 1;
assign key[877] = 648672;
assign key2[877] = 4753;
assign key3[877] = 1;
assign key[878] = 643921;
assign key2[878] = 4748;
assign key3[878] = 1;
assign key[879] = 639174;
assign key2[879] = 4743;
assign key3[879] = 1;
assign key[880] = 634433;
assign key2[880] = 4738;
assign key3[880] = 1;
assign key[881] = 629696;
assign key2[881] = 4734;
assign key3[881] = 1;
assign key[882] = 624965;
assign key2[882] = 4729;
assign key3[882] = 1;
assign key[883] = 620238;
assign key2[883] = 4724;
assign key3[883] = 1;
assign key[884] = 615517;
assign key2[884] = 4719;
assign key3[884] = 1;
assign key[885] = 610800;
assign key2[885] = 4714;
assign key3[885] = 1;
assign key[886] = 606088;
assign key2[886] = 4709;
assign key3[886] = 1;
assign key[887] = 601381;
assign key2[887] = 4704;
assign key3[887] = 1;
assign key[888] = 596680;
assign key2[888] = 4699;
assign key3[888] = 1;
assign key[889] = 591983;
assign key2[889] = 4694;
assign key3[889] = 1;
assign key[890] = 587291;
assign key2[890] = 4689;
assign key3[890] = 1;
assign key[891] = 582603;
assign key2[891] = 4684;
assign key3[891] = 1;
assign key[892] = 577921;
assign key2[892] = 4679;
assign key3[892] = 1;
assign key[893] = 573244;
assign key2[893] = 4674;
assign key3[893] = 1;
assign key[894] = 568571;
assign key2[894] = 4670;
assign key3[894] = 1;
assign key[895] = 563904;
assign key2[895] = 4665;
assign key3[895] = 1;
assign key[896] = 559241;
assign key2[896] = 4660;
assign key3[896] = 1;
assign key[897] = 554583;
assign key2[897] = 4655;
assign key3[897] = 1;
assign key[898] = 549930;
assign key2[898] = 4650;
assign key3[898] = 1;
assign key[899] = 545282;
assign key2[899] = 4645;
assign key3[899] = 1;
assign key[900] = 540638;
assign key2[900] = 4640;
assign key3[900] = 1;
assign key[901] = 536000;
assign key2[901] = 4636;
assign key3[901] = 1;
assign key[902] = 531366;
assign key2[902] = 4631;
assign key3[902] = 1;
assign key[903] = 526737;
assign key2[903] = 4626;
assign key3[903] = 1;
assign key[904] = 522113;
assign key2[904] = 4621;
assign key3[904] = 1;
assign key[905] = 517493;
assign key2[905] = 4616;
assign key3[905] = 1;
assign key[906] = 512879;
assign key2[906] = 4612;
assign key3[906] = 1;
assign key[907] = 508269;
assign key2[907] = 4607;
assign key3[907] = 1;
assign key[908] = 503664;
assign key2[908] = 4602;
assign key3[908] = 1;
assign key[909] = 499064;
assign key2[909] = 4597;
assign key3[909] = 1;
assign key[910] = 494468;
assign key2[910] = 4593;
assign key3[910] = 1;
assign key[911] = 489878;
assign key2[911] = 4588;
assign key3[911] = 1;
assign key[912] = 485292;
assign key2[912] = 4583;
assign key3[912] = 1;
assign key[913] = 480710;
assign key2[913] = 4578;
assign key3[913] = 1;
assign key[914] = 476134;
assign key2[914] = 4574;
assign key3[914] = 1;
assign key[915] = 471562;
assign key2[915] = 4569;
assign key3[915] = 1;
assign key[916] = 466995;
assign key2[916] = 4564;
assign key3[916] = 1;
assign key[917] = 462433;
assign key2[917] = 4560;
assign key3[917] = 1;
assign key[918] = 457875;
assign key2[918] = 4555;
assign key3[918] = 1;
assign key[919] = 453322;
assign key2[919] = 4550;
assign key3[919] = 1;
assign key[920] = 448774;
assign key2[920] = 4545;
assign key3[920] = 1;
assign key[921] = 444230;
assign key2[921] = 4541;
assign key3[921] = 1;
assign key[922] = 439691;
assign key2[922] = 4536;
assign key3[922] = 1;
assign key[923] = 435157;
assign key2[923] = 4531;
assign key3[923] = 1;
assign key[924] = 430627;
assign key2[924] = 4527;
assign key3[924] = 1;
assign key[925] = 426102;
assign key2[925] = 4522;
assign key3[925] = 1;
assign key[926] = 421582;
assign key2[926] = 4518;
assign key3[926] = 1;
assign key[927] = 417066;
assign key2[927] = 4513;
assign key3[927] = 1;
assign key[928] = 412555;
assign key2[928] = 4508;
assign key3[928] = 1;
assign key[929] = 408048;
assign key2[929] = 4504;
assign key3[929] = 1;
assign key[930] = 403546;
assign key2[930] = 4499;
assign key3[930] = 1;
assign key[931] = 399049;
assign key2[931] = 4494;
assign key3[931] = 1;
assign key[932] = 394556;
assign key2[932] = 4490;
assign key3[932] = 1;
assign key[933] = 390068;
assign key2[933] = 4485;
assign key3[933] = 1;
assign key[934] = 385585;
assign key2[934] = 4481;
assign key3[934] = 1;
assign key[935] = 381106;
assign key2[935] = 4476;
assign key3[935] = 1;
assign key[936] = 376632;
assign key2[936] = 4472;
assign key3[936] = 1;
assign key[937] = 372162;
assign key2[937] = 4467;
assign key3[937] = 1;
assign key[938] = 367697;
assign key2[938] = 4462;
assign key3[938] = 1;
assign key[939] = 363236;
assign key2[939] = 4458;
assign key3[939] = 1;
assign key[940] = 358780;
assign key2[940] = 4453;
assign key3[940] = 1;
assign key[941] = 354328;
assign key2[941] = 4449;
assign key3[941] = 1;
assign key[942] = 349881;
assign key2[942] = 4444;
assign key3[942] = 1;
assign key[943] = 345439;
assign key2[943] = 4440;
assign key3[943] = 1;
assign key[944] = 341001;
assign key2[944] = 4435;
assign key3[944] = 1;
assign key[945] = 336567;
assign key2[945] = 4431;
assign key3[945] = 1;
assign key[946] = 332138;
assign key2[946] = 4426;
assign key3[946] = 1;
assign key[947] = 327714;
assign key2[947] = 4422;
assign key3[947] = 1;
assign key[948] = 323293;
assign key2[948] = 4417;
assign key3[948] = 1;
assign key[949] = 318878;
assign key2[949] = 4413;
assign key3[949] = 1;
assign key[950] = 314467;
assign key2[950] = 4408;
assign key3[950] = 1;
assign key[951] = 310060;
assign key2[951] = 4404;
assign key3[951] = 1;
assign key[952] = 305658;
assign key2[952] = 4399;
assign key3[952] = 1;
assign key[953] = 301260;
assign key2[953] = 4395;
assign key3[953] = 1;
assign key[954] = 296867;
assign key2[954] = 4391;
assign key3[954] = 1;
assign key[955] = 292478;
assign key2[955] = 4386;
assign key3[955] = 1;
assign key[956] = 288094;
assign key2[956] = 4382;
assign key3[956] = 1;
assign key[957] = 283714;
assign key2[957] = 4377;
assign key3[957] = 1;
assign key[958] = 279338;
assign key2[958] = 4373;
assign key3[958] = 1;
assign key[959] = 274967;
assign key2[959] = 4368;
assign key3[959] = 1;
assign key[960] = 270601;
assign key2[960] = 4364;
assign key3[960] = 1;
assign key[961] = 266238;
assign key2[961] = 4360;
assign key3[961] = 1;
assign key[962] = 261880;
assign key2[962] = 4355;
assign key3[962] = 1;
assign key[963] = 257527;
assign key2[963] = 4351;
assign key3[963] = 1;
assign key[964] = 253178;
assign key2[964] = 4346;
assign key3[964] = 1;
assign key[965] = 248833;
assign key2[965] = 4342;
assign key3[965] = 1;
assign key[966] = 244492;
assign key2[966] = 4338;
assign key3[966] = 1;
assign key[967] = 240156;
assign key2[967] = 4333;
assign key3[967] = 1;
assign key[968] = 235825;
assign key2[968] = 4329;
assign key3[968] = 1;
assign key[969] = 231497;
assign key2[969] = 4325;
assign key3[969] = 1;
assign key[970] = 227174;
assign key2[970] = 4320;
assign key3[970] = 1;
assign key[971] = 222856;
assign key2[971] = 4316;
assign key3[971] = 1;
assign key[972] = 218541;
assign key2[972] = 4312;
assign key3[972] = 1;
assign key[973] = 214231;
assign key2[973] = 4307;
assign key3[973] = 1;
assign key[974] = 209925;
assign key2[974] = 4303;
assign key3[974] = 1;
assign key[975] = 205624;
assign key2[975] = 4299;
assign key3[975] = 1;
assign key[976] = 201327;
assign key2[976] = 4294;
assign key3[976] = 1;
assign key[977] = 197034;
assign key2[977] = 4290;
assign key3[977] = 1;
assign key[978] = 192746;
assign key2[978] = 4286;
assign key3[978] = 1;
assign key[979] = 188461;
assign key2[979] = 4282;
assign key3[979] = 1;
assign key[980] = 184181;
assign key2[980] = 4277;
assign key3[980] = 1;
assign key[981] = 179906;
assign key2[981] = 4273;
assign key3[981] = 1;
assign key[982] = 175634;
assign key2[982] = 4269;
assign key3[982] = 1;
assign key[983] = 171367;
assign key2[983] = 4265;
assign key3[983] = 1;
assign key[984] = 167104;
assign key2[984] = 4260;
assign key3[984] = 1;
assign key[985] = 162845;
assign key2[985] = 4256;
assign key3[985] = 1;
assign key[986] = 158591;
assign key2[986] = 4252;
assign key3[986] = 1;
assign key[987] = 154341;
assign key2[987] = 4248;
assign key3[987] = 1;
assign key[988] = 150095;
assign key2[988] = 4243;
assign key3[988] = 1;
assign key[989] = 145853;
assign key2[989] = 4239;
assign key3[989] = 1;
assign key[990] = 141615;
assign key2[990] = 4235;
assign key3[990] = 1;
assign key[991] = 137382;
assign key2[991] = 4231;
assign key3[991] = 1;
assign key[992] = 133153;
assign key2[992] = 4227;
assign key3[992] = 1;
assign key[993] = 128928;
assign key2[993] = 4222;
assign key3[993] = 1;
assign key[994] = 124707;
assign key2[994] = 4218;
assign key3[994] = 1;
assign key[995] = 120490;
assign key2[995] = 4214;
assign key3[995] = 1;
assign key[996] = 116278;
assign key2[996] = 4210;
assign key3[996] = 1;
assign key[997] = 112070;
assign key2[997] = 4206;
assign key3[997] = 1;
assign key[998] = 107866;
assign key2[998] = 4202;
assign key3[998] = 1;
assign key[999] = 103666;
assign key2[999] = 4197;
assign key3[999] = 1;
assign key[1000] = 99470;
assign key2[1000] = 4193;
assign key3[1000] = 1;
assign key[1001] = 95278;
assign key2[1001] = 4189;
assign key3[1001] = 1;
assign key[1002] = 91091;
assign key2[1002] = 4185;
assign key3[1002] = 1;
assign key[1003] = 86907;
assign key2[1003] = 4181;
assign key3[1003] = 1;
assign key[1004] = 82728;
assign key2[1004] = 4177;
assign key3[1004] = 1;
assign key[1005] = 78553;
assign key2[1005] = 4173;
assign key3[1005] = 1;
assign key[1006] = 74382;
assign key2[1006] = 4168;
assign key3[1006] = 1;
assign key[1007] = 70215;
assign key2[1007] = 4164;
assign key3[1007] = 1;
assign key[1008] = 66052;
assign key2[1008] = 4160;
assign key3[1008] = 1;
assign key[1009] = 61894;
assign key2[1009] = 4156;
assign key3[1009] = 1;
assign key[1010] = 57739;
assign key2[1010] = 4152;
assign key3[1010] = 1;
assign key[1011] = 53588;
assign key2[1011] = 4148;
assign key3[1011] = 1;
assign key[1012] = 49442;
assign key2[1012] = 4144;
assign key3[1012] = 1;
assign key[1013] = 45300;
assign key2[1013] = 4140;
assign key3[1013] = 1;
assign key[1014] = 41161;
assign key2[1014] = 4136;
assign key3[1014] = 1;
assign key[1015] = 37027;
assign key2[1015] = 4132;
assign key3[1015] = 1;
assign key[1016] = 32897;
assign key2[1016] = 4128;
assign key3[1016] = 1;
assign key[1017] = 28771;
assign key2[1017] = 4124;
assign key3[1017] = 1;
assign key[1018] = 24648;
assign key2[1018] = 4120;
assign key3[1018] = 1;
assign key[1019] = 20530;
assign key2[1019] = 4116;
assign key3[1019] = 1;
assign key[1020] = 16416;
assign key2[1020] = 4112;
assign key3[1020] = 1;
assign key[1021] = 12306;
assign key2[1021] = 4108;
assign key3[1021] = 1;
assign key[1022] = 8200;
assign key2[1022] = 4104;
assign key3[1022] = 1;
assign key[1023] = 4098;
assign key2[1023] = 4100;
assign key3[1023] = 1;
assign key[1024] = 0;
assign key2[1024] = 4096;
assign key3[1024] = 1;

wire [9:0] index;
assign index = bdata[22:13];

wire [22:0] a;
assign a = bdata[12] ? key[index+1] : key[index];

wire [12:0] b;
assign b = bdata[12:0];

wire [12:0] bb;
assign bb = ~bdata[12:0] + 1;

wire [25:0] bk;
assign bk = b * key2[index];

wire [25:0] bbk;
assign bbk = bb * key2[index+1];

wire c;
assign c = bdata[12] ? key3[index+1] : key3[index];

reg [22:0] a_reg;
reg [25:0] bk_reg;
reg [25:0] bbk_reg;
reg [31:0] adata_reg_1;
reg bs_reg_1;
reg [7:0] be_reg_1;
reg flag_reg_1;
reg [4:0] address_reg_1;
reg bdata12_reg;
reg c_reg;

always_ff@(posedge clk) begin
a_reg <= a;
bk_reg <= bk;
bbk_reg <= bbk;
adata_reg_1 <= adata;
bs_reg_1 <= bdata[31];
be_reg_1 <= bdata[30:23];
flag_reg_1 <= flag_in;
address_reg_1 <= address_in;
bdata12_reg <= bdata[12];
c_reg <= c;
end

wire [22:0] inv;
assign inv = bdata12_reg ? (c_reg ? a_reg + bbk_reg[25:13] : a_reg + bbk_reg[25:12]) : (c_reg ? a_reg - bk_reg[25:13] : a_reg - bk_reg[25:12]);

reg [31:0] adata_reg_2;
reg bs_reg_2;
reg [7:0] be_reg_2;
reg flag_reg_2;
reg [4:0] address_reg_2;
reg [22:0] inv_reg;

always_ff@(posedge clk) begin
adata_reg_2 <= adata_reg_1;
bs_reg_2 <= bs_reg_1;
be_reg_2 <= 253 - be_reg_1;
flag_reg_2 <= flag_reg_1;
address_reg_2 <= address_reg_1;
inv_reg <= inv;
end

wire [13:0] a0;
assign a0 = {1'b1,adata_reg_2[22:10]};

wire [13:0] b0;
assign b0 = {1'b1,inv_reg[22:10]};

wire [9:0] a1;
assign a1 = adata_reg_2[9:0];

wire [9:0] b1;
assign b1 = inv_reg[9:0];

wire [8:0] eadd;
assign eadd = adata_reg_2[30:23] + be_reg_2;

reg [27:0] a0b0;
reg [23:0] a1b0;
reg [23:0] a0b1;
reg [7:0] e;
reg [7:0] e_kuriage;
reg s;
reg notzero;
reg flag;
reg [4:0] address;

always@(posedge clk) begin

a0b0 <= a0 * b0;

a1b0 <= a1 * b0;

a0b1 <= a0 * b1;

e <= (eadd < 127) ? 0 : eadd - 127;

e_kuriage <= (eadd < 127) ? 0 : eadd - 126;

s <= adata_reg_2[31] ^ bs_reg_2;

notzero <= (|adata_reg_2[30:23]);

flag <= flag_reg_2;

address <= address_reg_2;

end

wire [14:0] a0b1tasua1b0;
assign a0b1tasua1b0 = a1b0[23:10] + a0b1[23:10] ;

wire [15:0] kekka_L;
assign kekka_L= a0b1tasua1b0 + a0b0[14:0];

wire [12:0] kekka_H_carry;
assign kekka_H_carry = a0b0[27:15] + 1;

wire [12:0] kekka_H_nocarry;
assign kekka_H_nocarry = a0b0[27:15];

wire carry;
assign carry = kekka_L[15];

wire [24:0] kekka;
assign kekka = carry ? {kekka_H_carry,kekka_L[14:3]} : {kekka_H_nocarry,kekka_L[14:3]};


wire [31:0] kotae;
assign kotae = notzero ? 
( kekka[24] ? {s,e_kuriage,kekka[23:1]} : {s,e,kekka[22:0]} ) : 0;

always@(posedge clk) begin
result <= kotae;
flag_out <= flag;
address_out <= address;
end
endmodule

`default_nettype wire


 


































