`default_nettype none

module fsqrt(
input wire [31:0] adata,
output reg [31:0] result,
input wire clk,
input wire flag_in,
input wire [4:0] address_in,
output reg flag_out,
output reg [4:0] address_out);

(* ram_style = "distributed" *) reg [22:0] s  [2047:0];
(* ram_style = "distributed" *) reg [12:0] tm [2047:0];
(* ram_style = "distributed" *) reg [5:0]  te [2047:0];

assign s[0] = 3474670;
assign tm[0] = 5796;
assign te[0] = 13;
assign s[1] = 3480462;
assign tm[1] = 5794;
assign te[1] = 13;
assign s[2] = 3486250;
assign tm[2] = 5791;
assign te[2] = 13;
assign s[3] = 3492035;
assign tm[3] = 5788;
assign te[3] = 13;
assign s[4] = 3497818;
assign tm[4] = 5785;
assign te[4] = 13;
assign s[5] = 3503598;
assign tm[5] = 5782;
assign te[5] = 13;
assign s[6] = 3509375;
assign tm[6] = 5779;
assign te[6] = 13;
assign s[7] = 3515149;
assign tm[7] = 5777;
assign te[7] = 13;
assign s[8] = 3520921;
assign tm[8] = 5774;
assign te[8] = 13;
assign s[9] = 3526689;
assign tm[9] = 5771;
assign te[9] = 13;
assign s[10] = 3532455;
assign tm[10] = 5768;
assign te[10] = 13;
assign s[11] = 3538218;
assign tm[11] = 5765;
assign te[11] = 13;
assign s[12] = 3543979;
assign tm[12] = 5763;
assign te[12] = 13;
assign s[13] = 3549737;
assign tm[13] = 5760;
assign te[13] = 13;
assign s[14] = 3555492;
assign tm[14] = 5757;
assign te[14] = 13;
assign s[15] = 3561244;
assign tm[15] = 5754;
assign te[15] = 13;
assign s[16] = 3566993;
assign tm[16] = 5752;
assign te[16] = 13;
assign s[17] = 3572739;
assign tm[17] = 5749;
assign te[17] = 13;
assign s[18] = 3578483;
assign tm[18] = 5746;
assign te[18] = 13;
assign s[19] = 3584224;
assign tm[19] = 5743;
assign te[19] = 13;
assign s[20] = 3589963;
assign tm[20] = 5740;
assign te[20] = 13;
assign s[21] = 3595698;
assign tm[21] = 5738;
assign te[21] = 13;
assign s[22] = 3601431;
assign tm[22] = 5735;
assign te[22] = 13;
assign s[23] = 3607160;
assign tm[23] = 5732;
assign te[23] = 13;
assign s[24] = 3612888;
assign tm[24] = 5730;
assign te[24] = 13;
assign s[25] = 3618613;
assign tm[25] = 5727;
assign te[25] = 13;
assign s[26] = 3624334;
assign tm[26] = 5724;
assign te[26] = 13;
assign s[27] = 3630053;
assign tm[27] = 5721;
assign te[27] = 13;
assign s[28] = 3635770;
assign tm[28] = 5719;
assign te[28] = 13;
assign s[29] = 3641484;
assign tm[29] = 5716;
assign te[29] = 13;
assign s[30] = 3647194;
assign tm[30] = 5713;
assign te[30] = 13;
assign s[31] = 3652903;
assign tm[31] = 5710;
assign te[31] = 13;
assign s[32] = 3658608;
assign tm[32] = 5708;
assign te[32] = 13;
assign s[33] = 3664311;
assign tm[33] = 5705;
assign te[33] = 13;
assign s[34] = 3670011;
assign tm[34] = 5702;
assign te[34] = 13;
assign s[35] = 3675708;
assign tm[35] = 5700;
assign te[35] = 13;
assign s[36] = 3681403;
assign tm[36] = 5697;
assign te[36] = 13;
assign s[37] = 3687095;
assign tm[37] = 5694;
assign te[37] = 13;
assign s[38] = 3692784;
assign tm[38] = 5692;
assign te[38] = 13;
assign s[39] = 3698471;
assign tm[39] = 5689;
assign te[39] = 13;
assign s[40] = 3704156;
assign tm[40] = 5686;
assign te[40] = 13;
assign s[41] = 3709837;
assign tm[41] = 5684;
assign te[41] = 13;
assign s[42] = 3715515;
assign tm[42] = 5681;
assign te[42] = 13;
assign s[43] = 3721191;
assign tm[43] = 5678;
assign te[43] = 13;
assign s[44] = 3726865;
assign tm[44] = 5676;
assign te[44] = 13;
assign s[45] = 3732536;
assign tm[45] = 5673;
assign te[45] = 13;
assign s[46] = 3738203;
assign tm[46] = 5670;
assign te[46] = 13;
assign s[47] = 3743869;
assign tm[47] = 5668;
assign te[47] = 13;
assign s[48] = 3749532;
assign tm[48] = 5665;
assign te[48] = 13;
assign s[49] = 3755192;
assign tm[49] = 5662;
assign te[49] = 13;
assign s[50] = 3760849;
assign tm[50] = 5660;
assign te[50] = 13;
assign s[51] = 3766504;
assign tm[51] = 5657;
assign te[51] = 13;
assign s[52] = 3772156;
assign tm[52] = 5654;
assign te[52] = 13;
assign s[53] = 3777806;
assign tm[53] = 5652;
assign te[53] = 13;
assign s[54] = 3783453;
assign tm[54] = 5649;
assign te[54] = 13;
assign s[55] = 3789097;
assign tm[55] = 5646;
assign te[55] = 13;
assign s[56] = 3794739;
assign tm[56] = 5644;
assign te[56] = 13;
assign s[57] = 3800378;
assign tm[57] = 5641;
assign te[57] = 13;
assign s[58] = 3806015;
assign tm[58] = 5639;
assign te[58] = 13;
assign s[59] = 3811648;
assign tm[59] = 5636;
assign te[59] = 13;
assign s[60] = 3817280;
assign tm[60] = 5633;
assign te[60] = 13;
assign s[61] = 3822909;
assign tm[61] = 5631;
assign te[61] = 13;
assign s[62] = 3828535;
assign tm[62] = 5628;
assign te[62] = 13;
assign s[63] = 3834158;
assign tm[63] = 5626;
assign te[63] = 13;
assign s[64] = 3839780;
assign tm[64] = 5623;
assign te[64] = 13;
assign s[65] = 3845398;
assign tm[65] = 5620;
assign te[65] = 13;
assign s[66] = 3851014;
assign tm[66] = 5618;
assign te[66] = 13;
assign s[67] = 3856626;
assign tm[67] = 5615;
assign te[67] = 13;
assign s[68] = 3862238;
assign tm[68] = 5613;
assign te[68] = 13;
assign s[69] = 3867846;
assign tm[69] = 5610;
assign te[69] = 13;
assign s[70] = 3873451;
assign tm[70] = 5608;
assign te[70] = 13;
assign s[71] = 3879054;
assign tm[71] = 5605;
assign te[71] = 13;
assign s[72] = 3884654;
assign tm[72] = 5602;
assign te[72] = 13;
assign s[73] = 3890253;
assign tm[73] = 5600;
assign te[73] = 13;
assign s[74] = 3895847;
assign tm[74] = 5597;
assign te[74] = 13;
assign s[75] = 3901440;
assign tm[75] = 5595;
assign te[75] = 13;
assign s[76] = 3907031;
assign tm[76] = 5592;
assign te[76] = 13;
assign s[77] = 3912618;
assign tm[77] = 5590;
assign te[77] = 13;
assign s[78] = 3918203;
assign tm[78] = 5587;
assign te[78] = 13;
assign s[79] = 3923786;
assign tm[79] = 5585;
assign te[79] = 13;
assign s[80] = 3929366;
assign tm[80] = 5582;
assign te[80] = 13;
assign s[81] = 3934944;
assign tm[81] = 5580;
assign te[81] = 13;
assign s[82] = 3940519;
assign tm[82] = 5577;
assign te[82] = 13;
assign s[83] = 3946091;
assign tm[83] = 5575;
assign te[83] = 13;
assign s[84] = 3951661;
assign tm[84] = 5572;
assign te[84] = 13;
assign s[85] = 3957229;
assign tm[85] = 5569;
assign te[85] = 13;
assign s[86] = 3962793;
assign tm[86] = 5567;
assign te[86] = 13;
assign s[87] = 3968356;
assign tm[87] = 5564;
assign te[87] = 13;
assign s[88] = 3973916;
assign tm[88] = 5562;
assign te[88] = 13;
assign s[89] = 3979474;
assign tm[89] = 5559;
assign te[89] = 13;
assign s[90] = 3985028;
assign tm[90] = 5557;
assign te[90] = 13;
assign s[91] = 3990581;
assign tm[91] = 5554;
assign te[91] = 13;
assign s[92] = 3996130;
assign tm[92] = 5552;
assign te[92] = 13;
assign s[93] = 4001678;
assign tm[93] = 5549;
assign te[93] = 13;
assign s[94] = 4007223;
assign tm[94] = 5547;
assign te[94] = 13;
assign s[95] = 4012766;
assign tm[95] = 5544;
assign te[95] = 13;
assign s[96] = 4018305;
assign tm[96] = 5542;
assign te[96] = 13;
assign s[97] = 4023843;
assign tm[97] = 5540;
assign te[97] = 13;
assign s[98] = 4029378;
assign tm[98] = 5537;
assign te[98] = 13;
assign s[99] = 4034911;
assign tm[99] = 5535;
assign te[99] = 13;
assign s[100] = 4040441;
assign tm[100] = 5532;
assign te[100] = 13;
assign s[101] = 4045969;
assign tm[101] = 5530;
assign te[101] = 13;
assign s[102] = 4051494;
assign tm[102] = 5527;
assign te[102] = 13;
assign s[103] = 4057017;
assign tm[103] = 5525;
assign te[103] = 13;
assign s[104] = 4062537;
assign tm[104] = 5522;
assign te[104] = 13;
assign s[105] = 4068055;
assign tm[105] = 5520;
assign te[105] = 13;
assign s[106] = 4073571;
assign tm[106] = 5517;
assign te[106] = 13;
assign s[107] = 4079084;
assign tm[107] = 5515;
assign te[107] = 13;
assign s[108] = 4084594;
assign tm[108] = 5513;
assign te[108] = 13;
assign s[109] = 4090102;
assign tm[109] = 5510;
assign te[109] = 13;
assign s[110] = 4095608;
assign tm[110] = 5508;
assign te[110] = 13;
assign s[111] = 4101112;
assign tm[111] = 5505;
assign te[111] = 13;
assign s[112] = 4106612;
assign tm[112] = 5503;
assign te[112] = 13;
assign s[113] = 4112111;
assign tm[113] = 5500;
assign te[113] = 13;
assign s[114] = 4117607;
assign tm[114] = 5498;
assign te[114] = 13;
assign s[115] = 4123100;
assign tm[115] = 5496;
assign te[115] = 13;
assign s[116] = 4128591;
assign tm[116] = 5493;
assign te[116] = 13;
assign s[117] = 4134080;
assign tm[117] = 5491;
assign te[117] = 13;
assign s[118] = 4139566;
assign tm[118] = 5488;
assign te[118] = 13;
assign s[119] = 4145050;
assign tm[119] = 5486;
assign te[119] = 13;
assign s[120] = 4150532;
assign tm[120] = 5483;
assign te[120] = 13;
assign s[121] = 4156011;
assign tm[121] = 5481;
assign te[121] = 13;
assign s[122] = 4161489;
assign tm[122] = 5479;
assign te[122] = 13;
assign s[123] = 4166963;
assign tm[123] = 5476;
assign te[123] = 13;
assign s[124] = 4172435;
assign tm[124] = 5474;
assign te[124] = 13;
assign s[125] = 4177904;
assign tm[125] = 5472;
assign te[125] = 13;
assign s[126] = 4183371;
assign tm[126] = 5469;
assign te[126] = 13;
assign s[127] = 4188837;
assign tm[127] = 5467;
assign te[127] = 13;
assign s[128] = 4194299;
assign tm[128] = 5464;
assign te[128] = 13;
assign s[129] = 4199760;
assign tm[129] = 5462;
assign te[129] = 13;
assign s[130] = 4205217;
assign tm[130] = 5460;
assign te[130] = 13;
assign s[131] = 4210673;
assign tm[131] = 5457;
assign te[131] = 13;
assign s[132] = 4216125;
assign tm[132] = 5455;
assign te[132] = 13;
assign s[133] = 4221577;
assign tm[133] = 5453;
assign te[133] = 13;
assign s[134] = 4227024;
assign tm[134] = 5450;
assign te[134] = 13;
assign s[135] = 4232470;
assign tm[135] = 5448;
assign te[135] = 13;
assign s[136] = 4237914;
assign tm[136] = 5445;
assign te[136] = 13;
assign s[137] = 4243355;
assign tm[137] = 5443;
assign te[137] = 13;
assign s[138] = 4248794;
assign tm[138] = 5441;
assign te[138] = 13;
assign s[139] = 4254231;
assign tm[139] = 5438;
assign te[139] = 13;
assign s[140] = 4259666;
assign tm[140] = 5436;
assign te[140] = 13;
assign s[141] = 4265097;
assign tm[141] = 5434;
assign te[141] = 13;
assign s[142] = 4270527;
assign tm[142] = 5431;
assign te[142] = 13;
assign s[143] = 4275954;
assign tm[143] = 5429;
assign te[143] = 13;
assign s[144] = 4281379;
assign tm[144] = 5427;
assign te[144] = 13;
assign s[145] = 4286801;
assign tm[145] = 5424;
assign te[145] = 13;
assign s[146] = 4292222;
assign tm[146] = 5422;
assign te[146] = 13;
assign s[147] = 4297640;
assign tm[147] = 5420;
assign te[147] = 13;
assign s[148] = 4303056;
assign tm[148] = 5417;
assign te[148] = 13;
assign s[149] = 4308470;
assign tm[149] = 5415;
assign te[149] = 13;
assign s[150] = 4313880;
assign tm[150] = 5413;
assign te[150] = 13;
assign s[151] = 4319289;
assign tm[151] = 5411;
assign te[151] = 13;
assign s[152] = 4324696;
assign tm[152] = 5408;
assign te[152] = 13;
assign s[153] = 4330100;
assign tm[153] = 5406;
assign te[153] = 13;
assign s[154] = 4335501;
assign tm[154] = 5404;
assign te[154] = 13;
assign s[155] = 4340901;
assign tm[155] = 5401;
assign te[155] = 13;
assign s[156] = 4346298;
assign tm[156] = 5399;
assign te[156] = 13;
assign s[157] = 4351694;
assign tm[157] = 5397;
assign te[157] = 13;
assign s[158] = 4357086;
assign tm[158] = 5394;
assign te[158] = 13;
assign s[159] = 4362477;
assign tm[159] = 5392;
assign te[159] = 13;
assign s[160] = 4367865;
assign tm[160] = 5390;
assign te[160] = 13;
assign s[161] = 4373251;
assign tm[161] = 5388;
assign te[161] = 13;
assign s[162] = 4378634;
assign tm[162] = 5385;
assign te[162] = 13;
assign s[163] = 4384016;
assign tm[163] = 5383;
assign te[163] = 13;
assign s[164] = 4389395;
assign tm[164] = 5381;
assign te[164] = 13;
assign s[165] = 4394772;
assign tm[165] = 5379;
assign te[165] = 13;
assign s[166] = 4400146;
assign tm[166] = 5376;
assign te[166] = 13;
assign s[167] = 4405519;
assign tm[167] = 5374;
assign te[167] = 13;
assign s[168] = 4410888;
assign tm[168] = 5372;
assign te[168] = 13;
assign s[169] = 4416257;
assign tm[169] = 5370;
assign te[169] = 13;
assign s[170] = 4421621;
assign tm[170] = 5367;
assign te[170] = 13;
assign s[171] = 4426985;
assign tm[171] = 5365;
assign te[171] = 13;
assign s[172] = 4432346;
assign tm[172] = 5363;
assign te[172] = 13;
assign s[173] = 4437705;
assign tm[173] = 5361;
assign te[173] = 13;
assign s[174] = 4443061;
assign tm[174] = 5358;
assign te[174] = 13;
assign s[175] = 4448416;
assign tm[175] = 5356;
assign te[175] = 13;
assign s[176] = 4453768;
assign tm[176] = 5354;
assign te[176] = 13;
assign s[177] = 4459118;
assign tm[177] = 5352;
assign te[177] = 13;
assign s[178] = 4464465;
assign tm[178] = 5349;
assign te[178] = 13;
assign s[179] = 4469811;
assign tm[179] = 5347;
assign te[179] = 13;
assign s[180] = 4475154;
assign tm[180] = 5345;
assign te[180] = 13;
assign s[181] = 4480495;
assign tm[181] = 5343;
assign te[181] = 13;
assign s[182] = 4485834;
assign tm[182] = 5340;
assign te[182] = 13;
assign s[183] = 4491170;
assign tm[183] = 5338;
assign te[183] = 13;
assign s[184] = 4496505;
assign tm[184] = 5336;
assign te[184] = 13;
assign s[185] = 4501837;
assign tm[185] = 5334;
assign te[185] = 13;
assign s[186] = 4507167;
assign tm[186] = 5332;
assign te[186] = 13;
assign s[187] = 4512494;
assign tm[187] = 5329;
assign te[187] = 13;
assign s[188] = 4517821;
assign tm[188] = 5327;
assign te[188] = 13;
assign s[189] = 4523144;
assign tm[189] = 5325;
assign te[189] = 13;
assign s[190] = 4528465;
assign tm[190] = 5323;
assign te[190] = 13;
assign s[191] = 4533783;
assign tm[191] = 5321;
assign te[191] = 13;
assign s[192] = 4539100;
assign tm[192] = 5318;
assign te[192] = 13;
assign s[193] = 4544415;
assign tm[193] = 5316;
assign te[193] = 13;
assign s[194] = 4549727;
assign tm[194] = 5314;
assign te[194] = 13;
assign s[195] = 4555038;
assign tm[195] = 5312;
assign te[195] = 13;
assign s[196] = 4560346;
assign tm[196] = 5310;
assign te[196] = 13;
assign s[197] = 4565651;
assign tm[197] = 5308;
assign te[197] = 13;
assign s[198] = 4570955;
assign tm[198] = 5305;
assign te[198] = 13;
assign s[199] = 4576257;
assign tm[199] = 5303;
assign te[199] = 13;
assign s[200] = 4581555;
assign tm[200] = 5301;
assign te[200] = 13;
assign s[201] = 4586853;
assign tm[201] = 5299;
assign te[201] = 13;
assign s[202] = 4592149;
assign tm[202] = 5297;
assign te[202] = 13;
assign s[203] = 4597441;
assign tm[203] = 5295;
assign te[203] = 13;
assign s[204] = 4602732;
assign tm[204] = 5292;
assign te[204] = 13;
assign s[205] = 4608020;
assign tm[205] = 5290;
assign te[205] = 13;
assign s[206] = 4613307;
assign tm[206] = 5288;
assign te[206] = 13;
assign s[207] = 4618591;
assign tm[207] = 5286;
assign te[207] = 13;
assign s[208] = 4623873;
assign tm[208] = 5284;
assign te[208] = 13;
assign s[209] = 4629153;
assign tm[209] = 5282;
assign te[209] = 13;
assign s[210] = 4634431;
assign tm[210] = 5279;
assign te[210] = 13;
assign s[211] = 4639706;
assign tm[211] = 5277;
assign te[211] = 13;
assign s[212] = 4644980;
assign tm[212] = 5275;
assign te[212] = 13;
assign s[213] = 4650252;
assign tm[213] = 5273;
assign te[213] = 13;
assign s[214] = 4655520;
assign tm[214] = 5271;
assign te[214] = 13;
assign s[215] = 4660788;
assign tm[215] = 5269;
assign te[215] = 13;
assign s[216] = 4666053;
assign tm[216] = 5267;
assign te[216] = 13;
assign s[217] = 4671316;
assign tm[217] = 5265;
assign te[217] = 13;
assign s[218] = 4676578;
assign tm[218] = 5262;
assign te[218] = 13;
assign s[219] = 4681836;
assign tm[219] = 5260;
assign te[219] = 13;
assign s[220] = 4687092;
assign tm[220] = 5258;
assign te[220] = 13;
assign s[221] = 4692346;
assign tm[221] = 5256;
assign te[221] = 13;
assign s[222] = 4697599;
assign tm[222] = 5254;
assign te[222] = 13;
assign s[223] = 4702849;
assign tm[223] = 5252;
assign te[223] = 13;
assign s[224] = 4708097;
assign tm[224] = 5250;
assign te[224] = 13;
assign s[225] = 4713344;
assign tm[225] = 5248;
assign te[225] = 13;
assign s[226] = 4718587;
assign tm[226] = 5246;
assign te[226] = 13;
assign s[227] = 4723829;
assign tm[227] = 5243;
assign te[227] = 13;
assign s[228] = 4729069;
assign tm[228] = 5241;
assign te[228] = 13;
assign s[229] = 4734306;
assign tm[229] = 5239;
assign te[229] = 13;
assign s[230] = 4739542;
assign tm[230] = 5237;
assign te[230] = 13;
assign s[231] = 4744776;
assign tm[231] = 5235;
assign te[231] = 13;
assign s[232] = 4750007;
assign tm[232] = 5233;
assign te[232] = 13;
assign s[233] = 4755236;
assign tm[233] = 5231;
assign te[233] = 13;
assign s[234] = 4760463;
assign tm[234] = 5229;
assign te[234] = 13;
assign s[235] = 4765689;
assign tm[235] = 5227;
assign te[235] = 13;
assign s[236] = 4770912;
assign tm[236] = 5225;
assign te[236] = 13;
assign s[237] = 4776133;
assign tm[237] = 5223;
assign te[237] = 13;
assign s[238] = 4781351;
assign tm[238] = 5220;
assign te[238] = 13;
assign s[239] = 4786569;
assign tm[239] = 5218;
assign te[239] = 13;
assign s[240] = 4791783;
assign tm[240] = 5216;
assign te[240] = 13;
assign s[241] = 4796996;
assign tm[241] = 5214;
assign te[241] = 13;
assign s[242] = 4802207;
assign tm[242] = 5212;
assign te[242] = 13;
assign s[243] = 4807416;
assign tm[243] = 5210;
assign te[243] = 13;
assign s[244] = 4812622;
assign tm[244] = 5208;
assign te[244] = 13;
assign s[245] = 4817827;
assign tm[245] = 5206;
assign te[245] = 13;
assign s[246] = 4823029;
assign tm[246] = 5204;
assign te[246] = 13;
assign s[247] = 4828230;
assign tm[247] = 5202;
assign te[247] = 13;
assign s[248] = 4833427;
assign tm[248] = 5200;
assign te[248] = 13;
assign s[249] = 4838624;
assign tm[249] = 5198;
assign te[249] = 13;
assign s[250] = 4843818;
assign tm[250] = 5196;
assign te[250] = 13;
assign s[251] = 4849010;
assign tm[251] = 5194;
assign te[251] = 13;
assign s[252] = 4854201;
assign tm[252] = 5192;
assign te[252] = 13;
assign s[253] = 4859389;
assign tm[253] = 5190;
assign te[253] = 13;
assign s[254] = 4864575;
assign tm[254] = 5188;
assign te[254] = 13;
assign s[255] = 4869759;
assign tm[255] = 5186;
assign te[255] = 13;
assign s[256] = 4874941;
assign tm[256] = 5184;
assign te[256] = 13;
assign s[257] = 4880121;
assign tm[257] = 5182;
assign te[257] = 13;
assign s[258] = 4885300;
assign tm[258] = 5180;
assign te[258] = 13;
assign s[259] = 4890475;
assign tm[259] = 5178;
assign te[259] = 13;
assign s[260] = 4895649;
assign tm[260] = 5176;
assign te[260] = 13;
assign s[261] = 4900821;
assign tm[261] = 5174;
assign te[261] = 13;
assign s[262] = 4905990;
assign tm[262] = 5171;
assign te[262] = 13;
assign s[263] = 4911159;
assign tm[263] = 5169;
assign te[263] = 13;
assign s[264] = 4916325;
assign tm[264] = 5167;
assign te[264] = 13;
assign s[265] = 4921489;
assign tm[265] = 5165;
assign te[265] = 13;
assign s[266] = 4926651;
assign tm[266] = 5163;
assign te[266] = 13;
assign s[267] = 4931811;
assign tm[267] = 5161;
assign te[267] = 13;
assign s[268] = 4936969;
assign tm[268] = 5159;
assign te[268] = 13;
assign s[269] = 4942124;
assign tm[269] = 5157;
assign te[269] = 13;
assign s[270] = 4947279;
assign tm[270] = 5155;
assign te[270] = 13;
assign s[271] = 4952431;
assign tm[271] = 5153;
assign te[271] = 13;
assign s[272] = 4957581;
assign tm[272] = 5151;
assign te[272] = 13;
assign s[273] = 4962729;
assign tm[273] = 5149;
assign te[273] = 13;
assign s[274] = 4967874;
assign tm[274] = 5147;
assign te[274] = 13;
assign s[275] = 4973019;
assign tm[275] = 5146;
assign te[275] = 13;
assign s[276] = 4978161;
assign tm[276] = 5144;
assign te[276] = 13;
assign s[277] = 4983301;
assign tm[277] = 5142;
assign te[277] = 13;
assign s[278] = 4988439;
assign tm[278] = 5140;
assign te[278] = 13;
assign s[279] = 4993576;
assign tm[279] = 5138;
assign te[279] = 13;
assign s[280] = 4998710;
assign tm[280] = 5136;
assign te[280] = 13;
assign s[281] = 5003842;
assign tm[281] = 5134;
assign te[281] = 13;
assign s[282] = 5008972;
assign tm[282] = 5132;
assign te[282] = 13;
assign s[283] = 5014100;
assign tm[283] = 5130;
assign te[283] = 13;
assign s[284] = 5019227;
assign tm[284] = 5128;
assign te[284] = 13;
assign s[285] = 5024351;
assign tm[285] = 5126;
assign te[285] = 13;
assign s[286] = 5029473;
assign tm[286] = 5124;
assign te[286] = 13;
assign s[287] = 5034593;
assign tm[287] = 5122;
assign te[287] = 13;
assign s[288] = 5039712;
assign tm[288] = 5120;
assign te[288] = 13;
assign s[289] = 5044828;
assign tm[289] = 5118;
assign te[289] = 13;
assign s[290] = 5049943;
assign tm[290] = 5116;
assign te[290] = 13;
assign s[291] = 5055056;
assign tm[291] = 5114;
assign te[291] = 13;
assign s[292] = 5060166;
assign tm[292] = 5112;
assign te[292] = 13;
assign s[293] = 5065275;
assign tm[293] = 5110;
assign te[293] = 13;
assign s[294] = 5070383;
assign tm[294] = 5108;
assign te[294] = 13;
assign s[295] = 5075487;
assign tm[295] = 5106;
assign te[295] = 13;
assign s[296] = 5080590;
assign tm[296] = 5104;
assign te[296] = 13;
assign s[297] = 5085691;
assign tm[297] = 5102;
assign te[297] = 13;
assign s[298] = 5090790;
assign tm[298] = 5101;
assign te[298] = 13;
assign s[299] = 5095887;
assign tm[299] = 5099;
assign te[299] = 13;
assign s[300] = 5100982;
assign tm[300] = 5097;
assign te[300] = 13;
assign s[301] = 5106076;
assign tm[301] = 5095;
assign te[301] = 13;
assign s[302] = 5111167;
assign tm[302] = 5093;
assign te[302] = 13;
assign s[303] = 5116257;
assign tm[303] = 5091;
assign te[303] = 13;
assign s[304] = 5121344;
assign tm[304] = 5089;
assign te[304] = 13;
assign s[305] = 5126430;
assign tm[305] = 5087;
assign te[305] = 13;
assign s[306] = 5131513;
assign tm[306] = 5085;
assign te[306] = 13;
assign s[307] = 5136595;
assign tm[307] = 5083;
assign te[307] = 13;
assign s[308] = 5141675;
assign tm[308] = 5081;
assign te[308] = 13;
assign s[309] = 5146753;
assign tm[309] = 5079;
assign te[309] = 13;
assign s[310] = 5151829;
assign tm[310] = 5077;
assign te[310] = 13;
assign s[311] = 5156903;
assign tm[311] = 5076;
assign te[311] = 13;
assign s[312] = 5161976;
assign tm[312] = 5074;
assign te[312] = 13;
assign s[313] = 5167046;
assign tm[313] = 5072;
assign te[313] = 13;
assign s[314] = 5172115;
assign tm[314] = 5070;
assign te[314] = 13;
assign s[315] = 5177181;
assign tm[315] = 5068;
assign te[315] = 13;
assign s[316] = 5182246;
assign tm[316] = 5066;
assign te[316] = 13;
assign s[317] = 5187308;
assign tm[317] = 5064;
assign te[317] = 13;
assign s[318] = 5192369;
assign tm[318] = 5062;
assign te[318] = 13;
assign s[319] = 5197428;
assign tm[319] = 5060;
assign te[319] = 13;
assign s[320] = 5202486;
assign tm[320] = 5059;
assign te[320] = 13;
assign s[321] = 5207541;
assign tm[321] = 5057;
assign te[321] = 13;
assign s[322] = 5212594;
assign tm[322] = 5055;
assign te[322] = 13;
assign s[323] = 5217646;
assign tm[323] = 5053;
assign te[323] = 13;
assign s[324] = 5222696;
assign tm[324] = 5051;
assign te[324] = 13;
assign s[325] = 5227744;
assign tm[325] = 5049;
assign te[325] = 13;
assign s[326] = 5232789;
assign tm[326] = 5047;
assign te[326] = 13;
assign s[327] = 5237833;
assign tm[327] = 5045;
assign te[327] = 13;
assign s[328] = 5242875;
assign tm[328] = 5044;
assign te[328] = 13;
assign s[329] = 5247916;
assign tm[329] = 5042;
assign te[329] = 13;
assign s[330] = 5252954;
assign tm[330] = 5040;
assign te[330] = 13;
assign s[331] = 5257991;
assign tm[331] = 5038;
assign te[331] = 13;
assign s[332] = 5263025;
assign tm[332] = 5036;
assign te[332] = 13;
assign s[333] = 5268058;
assign tm[333] = 5034;
assign te[333] = 13;
assign s[334] = 5273089;
assign tm[334] = 5032;
assign te[334] = 13;
assign s[335] = 5278118;
assign tm[335] = 5031;
assign te[335] = 13;
assign s[336] = 5283145;
assign tm[336] = 5029;
assign te[336] = 13;
assign s[337] = 5288172;
assign tm[337] = 5027;
assign te[337] = 13;
assign s[338] = 5293195;
assign tm[338] = 5025;
assign te[338] = 13;
assign s[339] = 5298216;
assign tm[339] = 5023;
assign te[339] = 13;
assign s[340] = 5303237;
assign tm[340] = 5021;
assign te[340] = 13;
assign s[341] = 5308255;
assign tm[341] = 5019;
assign te[341] = 13;
assign s[342] = 5313271;
assign tm[342] = 5018;
assign te[342] = 13;
assign s[343] = 5318285;
assign tm[343] = 5016;
assign te[343] = 13;
assign s[344] = 5323297;
assign tm[344] = 5014;
assign te[344] = 13;
assign s[345] = 5328308;
assign tm[345] = 5012;
assign te[345] = 13;
assign s[346] = 5333318;
assign tm[346] = 5010;
assign te[346] = 13;
assign s[347] = 5338324;
assign tm[347] = 5008;
assign te[347] = 13;
assign s[348] = 5343330;
assign tm[348] = 5007;
assign te[348] = 13;
assign s[349] = 5348333;
assign tm[349] = 5005;
assign te[349] = 13;
assign s[350] = 5353335;
assign tm[350] = 5003;
assign te[350] = 13;
assign s[351] = 5358334;
assign tm[351] = 5001;
assign te[351] = 13;
assign s[352] = 5363333;
assign tm[352] = 4999;
assign te[352] = 13;
assign s[353] = 5368329;
assign tm[353] = 4997;
assign te[353] = 13;
assign s[354] = 5373324;
assign tm[354] = 4996;
assign te[354] = 13;
assign s[355] = 5378315;
assign tm[355] = 4994;
assign te[355] = 13;
assign s[356] = 5383306;
assign tm[356] = 4992;
assign te[356] = 13;
assign s[357] = 5388295;
assign tm[357] = 4990;
assign te[357] = 13;
assign s[358] = 5393283;
assign tm[358] = 4988;
assign te[358] = 13;
assign s[359] = 5398268;
assign tm[359] = 4987;
assign te[359] = 13;
assign s[360] = 5403251;
assign tm[360] = 4985;
assign te[360] = 13;
assign s[361] = 5408233;
assign tm[361] = 4983;
assign te[361] = 13;
assign s[362] = 5413213;
assign tm[362] = 4981;
assign te[362] = 13;
assign s[363] = 5418191;
assign tm[363] = 4979;
assign te[363] = 13;
assign s[364] = 5423167;
assign tm[364] = 4978;
assign te[364] = 13;
assign s[365] = 5428142;
assign tm[365] = 4976;
assign te[365] = 13;
assign s[366] = 5433115;
assign tm[366] = 4974;
assign te[366] = 13;
assign s[367] = 5438086;
assign tm[367] = 4972;
assign te[367] = 13;
assign s[368] = 5443054;
assign tm[368] = 4970;
assign te[368] = 13;
assign s[369] = 5448023;
assign tm[369] = 4969;
assign te[369] = 13;
assign s[370] = 5452988;
assign tm[370] = 4967;
assign te[370] = 13;
assign s[371] = 5457952;
assign tm[371] = 4965;
assign te[371] = 13;
assign s[372] = 5462914;
assign tm[372] = 4963;
assign te[372] = 13;
assign s[373] = 5467874;
assign tm[373] = 4962;
assign te[373] = 13;
assign s[374] = 5472833;
assign tm[374] = 4960;
assign te[374] = 13;
assign s[375] = 5477789;
assign tm[375] = 4958;
assign te[375] = 13;
assign s[376] = 5482744;
assign tm[376] = 4956;
assign te[376] = 13;
assign s[377] = 5487697;
assign tm[377] = 4954;
assign te[377] = 13;
assign s[378] = 5492649;
assign tm[378] = 4953;
assign te[378] = 13;
assign s[379] = 5497598;
assign tm[379] = 4951;
assign te[379] = 13;
assign s[380] = 5502546;
assign tm[380] = 4949;
assign te[380] = 13;
assign s[381] = 5507493;
assign tm[381] = 4947;
assign te[381] = 13;
assign s[382] = 5512437;
assign tm[382] = 4946;
assign te[382] = 13;
assign s[383] = 5517379;
assign tm[383] = 4944;
assign te[383] = 13;
assign s[384] = 5522320;
assign tm[384] = 4942;
assign te[384] = 13;
assign s[385] = 5527259;
assign tm[385] = 4940;
assign te[385] = 13;
assign s[386] = 5532196;
assign tm[386] = 4939;
assign te[386] = 13;
assign s[387] = 5537132;
assign tm[387] = 4937;
assign te[387] = 13;
assign s[388] = 5542066;
assign tm[388] = 4935;
assign te[388] = 13;
assign s[389] = 5546998;
assign tm[389] = 4933;
assign te[389] = 13;
assign s[390] = 5551928;
assign tm[390] = 4932;
assign te[390] = 13;
assign s[391] = 5556857;
assign tm[391] = 4930;
assign te[391] = 13;
assign s[392] = 5561784;
assign tm[392] = 4928;
assign te[392] = 13;
assign s[393] = 5566709;
assign tm[393] = 4926;
assign te[393] = 13;
assign s[394] = 5571633;
assign tm[394] = 4925;
assign te[394] = 13;
assign s[395] = 5576554;
assign tm[395] = 4923;
assign te[395] = 13;
assign s[396] = 5581474;
assign tm[396] = 4921;
assign te[396] = 13;
assign s[397] = 5586392;
assign tm[397] = 4919;
assign te[397] = 13;
assign s[398] = 5591308;
assign tm[398] = 4918;
assign te[398] = 13;
assign s[399] = 5596223;
assign tm[399] = 4916;
assign te[399] = 13;
assign s[400] = 5601137;
assign tm[400] = 4914;
assign te[400] = 13;
assign s[401] = 5606047;
assign tm[401] = 4912;
assign te[401] = 13;
assign s[402] = 5610957;
assign tm[402] = 4911;
assign te[402] = 13;
assign s[403] = 5615865;
assign tm[403] = 4909;
assign te[403] = 13;
assign s[404] = 5620771;
assign tm[404] = 4907;
assign te[404] = 13;
assign s[405] = 5625675;
assign tm[405] = 4906;
assign te[405] = 13;
assign s[406] = 5630577;
assign tm[406] = 4904;
assign te[406] = 13;
assign s[407] = 5635478;
assign tm[407] = 4902;
assign te[407] = 13;
assign s[408] = 5640378;
assign tm[408] = 4900;
assign te[408] = 13;
assign s[409] = 5645275;
assign tm[409] = 4899;
assign te[409] = 13;
assign s[410] = 5650172;
assign tm[410] = 4897;
assign te[410] = 13;
assign s[411] = 5655066;
assign tm[411] = 4895;
assign te[411] = 13;
assign s[412] = 5659958;
assign tm[412] = 4894;
assign te[412] = 13;
assign s[413] = 5664849;
assign tm[413] = 4892;
assign te[413] = 13;
assign s[414] = 5669737;
assign tm[414] = 4890;
assign te[414] = 13;
assign s[415] = 5674625;
assign tm[415] = 4889;
assign te[415] = 13;
assign s[416] = 5679510;
assign tm[416] = 4887;
assign te[416] = 13;
assign s[417] = 5684395;
assign tm[417] = 4885;
assign te[417] = 13;
assign s[418] = 5689276;
assign tm[418] = 4883;
assign te[418] = 13;
assign s[419] = 5694157;
assign tm[419] = 4882;
assign te[419] = 13;
assign s[420] = 5699036;
assign tm[420] = 4880;
assign te[420] = 13;
assign s[421] = 5703914;
assign tm[421] = 4878;
assign te[421] = 13;
assign s[422] = 5708789;
assign tm[422] = 4877;
assign te[422] = 13;
assign s[423] = 5713663;
assign tm[423] = 4875;
assign te[423] = 13;
assign s[424] = 5718535;
assign tm[424] = 4873;
assign te[424] = 13;
assign s[425] = 5723405;
assign tm[425] = 4872;
assign te[425] = 13;
assign s[426] = 5728274;
assign tm[426] = 4870;
assign te[426] = 13;
assign s[427] = 5733141;
assign tm[427] = 4868;
assign te[427] = 13;
assign s[428] = 5738006;
assign tm[428] = 4867;
assign te[428] = 13;
assign s[429] = 5742870;
assign tm[429] = 4865;
assign te[429] = 13;
assign s[430] = 5747732;
assign tm[430] = 4863;
assign te[430] = 13;
assign s[431] = 5752593;
assign tm[431] = 4862;
assign te[431] = 13;
assign s[432] = 5757451;
assign tm[432] = 4860;
assign te[432] = 13;
assign s[433] = 5762308;
assign tm[433] = 4858;
assign te[433] = 13;
assign s[434] = 5767163;
assign tm[434] = 4857;
assign te[434] = 13;
assign s[435] = 5772017;
assign tm[435] = 4855;
assign te[435] = 13;
assign s[436] = 5776869;
assign tm[436] = 4853;
assign te[436] = 13;
assign s[437] = 5781719;
assign tm[437] = 4852;
assign te[437] = 13;
assign s[438] = 5786568;
assign tm[438] = 4850;
assign te[438] = 13;
assign s[439] = 5791416;
assign tm[439] = 4848;
assign te[439] = 13;
assign s[440] = 5796261;
assign tm[440] = 4847;
assign te[440] = 13;
assign s[441] = 5801105;
assign tm[441] = 4845;
assign te[441] = 13;
assign s[442] = 5805947;
assign tm[442] = 4843;
assign te[442] = 13;
assign s[443] = 5810787;
assign tm[443] = 4842;
assign te[443] = 13;
assign s[444] = 5815626;
assign tm[444] = 4840;
assign te[444] = 13;
assign s[445] = 5820463;
assign tm[445] = 4838;
assign te[445] = 13;
assign s[446] = 5825298;
assign tm[446] = 4837;
assign te[446] = 13;
assign s[447] = 5830132;
assign tm[447] = 4835;
assign te[447] = 13;
assign s[448] = 5834964;
assign tm[448] = 4833;
assign te[448] = 13;
assign s[449] = 5839795;
assign tm[449] = 4832;
assign te[449] = 13;
assign s[450] = 5844624;
assign tm[450] = 4830;
assign te[450] = 13;
assign s[451] = 5849451;
assign tm[451] = 4828;
assign te[451] = 13;
assign s[452] = 5854277;
assign tm[452] = 4827;
assign te[452] = 13;
assign s[453] = 5859100;
assign tm[453] = 4825;
assign te[453] = 13;
assign s[454] = 5863923;
assign tm[454] = 4824;
assign te[454] = 13;
assign s[455] = 5868744;
assign tm[455] = 4822;
assign te[455] = 13;
assign s[456] = 5873563;
assign tm[456] = 4820;
assign te[456] = 13;
assign s[457] = 5878380;
assign tm[457] = 4819;
assign te[457] = 13;
assign s[458] = 5883196;
assign tm[458] = 4817;
assign te[458] = 13;
assign s[459] = 5888010;
assign tm[459] = 4815;
assign te[459] = 13;
assign s[460] = 5892823;
assign tm[460] = 4814;
assign te[460] = 13;
assign s[461] = 5897634;
assign tm[461] = 4812;
assign te[461] = 13;
assign s[462] = 5902443;
assign tm[462] = 4810;
assign te[462] = 13;
assign s[463] = 5907251;
assign tm[463] = 4809;
assign te[463] = 13;
assign s[464] = 5912057;
assign tm[464] = 4807;
assign te[464] = 13;
assign s[465] = 5916862;
assign tm[465] = 4806;
assign te[465] = 13;
assign s[466] = 5921664;
assign tm[466] = 4804;
assign te[466] = 13;
assign s[467] = 5926466;
assign tm[467] = 4802;
assign te[467] = 13;
assign s[468] = 5931266;
assign tm[468] = 4801;
assign te[468] = 13;
assign s[469] = 5936064;
assign tm[469] = 4799;
assign te[469] = 13;
assign s[470] = 5940860;
assign tm[470] = 4798;
assign te[470] = 13;
assign s[471] = 5945656;
assign tm[471] = 4796;
assign te[471] = 13;
assign s[472] = 5950449;
assign tm[472] = 4794;
assign te[472] = 13;
assign s[473] = 5955240;
assign tm[473] = 4793;
assign te[473] = 13;
assign s[474] = 5960030;
assign tm[474] = 4791;
assign te[474] = 13;
assign s[475] = 5964819;
assign tm[475] = 4790;
assign te[475] = 13;
assign s[476] = 5969606;
assign tm[476] = 4788;
assign te[476] = 13;
assign s[477] = 5974391;
assign tm[477] = 4786;
assign te[477] = 13;
assign s[478] = 5979175;
assign tm[478] = 4785;
assign te[478] = 13;
assign s[479] = 5983957;
assign tm[479] = 4783;
assign te[479] = 13;
assign s[480] = 5988737;
assign tm[480] = 4782;
assign te[480] = 13;
assign s[481] = 5993517;
assign tm[481] = 4780;
assign te[481] = 13;
assign s[482] = 5998293;
assign tm[482] = 4778;
assign te[482] = 13;
assign s[483] = 6003069;
assign tm[483] = 4777;
assign te[483] = 13;
assign s[484] = 6007844;
assign tm[484] = 4775;
assign te[484] = 13;
assign s[485] = 6012616;
assign tm[485] = 4774;
assign te[485] = 13;
assign s[486] = 6017387;
assign tm[486] = 4772;
assign te[486] = 13;
assign s[487] = 6022157;
assign tm[487] = 4770;
assign te[487] = 13;
assign s[488] = 6026924;
assign tm[488] = 4769;
assign te[488] = 13;
assign s[489] = 6031691;
assign tm[489] = 4767;
assign te[489] = 13;
assign s[490] = 6036455;
assign tm[490] = 4766;
assign te[490] = 13;
assign s[491] = 6041219;
assign tm[491] = 4764;
assign te[491] = 13;
assign s[492] = 6045980;
assign tm[492] = 4763;
assign te[492] = 13;
assign s[493] = 6050740;
assign tm[493] = 4761;
assign te[493] = 13;
assign s[494] = 6055498;
assign tm[494] = 4759;
assign te[494] = 13;
assign s[495] = 6060255;
assign tm[495] = 4758;
assign te[495] = 13;
assign s[496] = 6065010;
assign tm[496] = 4756;
assign te[496] = 13;
assign s[497] = 6069764;
assign tm[497] = 4755;
assign te[497] = 13;
assign s[498] = 6074515;
assign tm[498] = 4753;
assign te[498] = 13;
assign s[499] = 6079267;
assign tm[499] = 4752;
assign te[499] = 13;
assign s[500] = 6084015;
assign tm[500] = 4750;
assign te[500] = 13;
assign s[501] = 6088763;
assign tm[501] = 4749;
assign te[501] = 13;
assign s[502] = 6093510;
assign tm[502] = 4747;
assign te[502] = 13;
assign s[503] = 6098253;
assign tm[503] = 4745;
assign te[503] = 13;
assign s[504] = 6102996;
assign tm[504] = 4744;
assign te[504] = 13;
assign s[505] = 6107737;
assign tm[505] = 4742;
assign te[505] = 13;
assign s[506] = 6112477;
assign tm[506] = 4741;
assign te[506] = 13;
assign s[507] = 6117215;
assign tm[507] = 4739;
assign te[507] = 13;
assign s[508] = 6121952;
assign tm[508] = 4738;
assign te[508] = 13;
assign s[509] = 6126687;
assign tm[509] = 4736;
assign te[509] = 13;
assign s[510] = 6131421;
assign tm[510] = 4735;
assign te[510] = 13;
assign s[511] = 6136152;
assign tm[511] = 4733;
assign te[511] = 13;
assign s[512] = 6140883;
assign tm[512] = 4731;
assign te[512] = 13;
assign s[513] = 6145611;
assign tm[513] = 4730;
assign te[513] = 13;
assign s[514] = 6150339;
assign tm[514] = 4728;
assign te[514] = 13;
assign s[515] = 6155065;
assign tm[515] = 4727;
assign te[515] = 13;
assign s[516] = 6159789;
assign tm[516] = 4725;
assign te[516] = 13;
assign s[517] = 6164511;
assign tm[517] = 4724;
assign te[517] = 13;
assign s[518] = 6169233;
assign tm[518] = 4722;
assign te[518] = 13;
assign s[519] = 6173953;
assign tm[519] = 4721;
assign te[519] = 13;
assign s[520] = 6178670;
assign tm[520] = 4719;
assign te[520] = 13;
assign s[521] = 6183388;
assign tm[521] = 4718;
assign te[521] = 13;
assign s[522] = 6188103;
assign tm[522] = 4716;
assign te[522] = 13;
assign s[523] = 6192816;
assign tm[523] = 4715;
assign te[523] = 13;
assign s[524] = 6197528;
assign tm[524] = 4713;
assign te[524] = 13;
assign s[525] = 6202239;
assign tm[525] = 4712;
assign te[525] = 13;
assign s[526] = 6206948;
assign tm[526] = 4710;
assign te[526] = 13;
assign s[527] = 6211655;
assign tm[527] = 4709;
assign te[527] = 13;
assign s[528] = 6216361;
assign tm[528] = 4707;
assign te[528] = 13;
assign s[529] = 6221066;
assign tm[529] = 4705;
assign te[529] = 13;
assign s[530] = 6225769;
assign tm[530] = 4704;
assign te[530] = 13;
assign s[531] = 6230470;
assign tm[531] = 4702;
assign te[531] = 13;
assign s[532] = 6235170;
assign tm[532] = 4701;
assign te[532] = 13;
assign s[533] = 6239868;
assign tm[533] = 4699;
assign te[533] = 13;
assign s[534] = 6244565;
assign tm[534] = 4698;
assign te[534] = 13;
assign s[535] = 6249261;
assign tm[535] = 4696;
assign te[535] = 13;
assign s[536] = 6253954;
assign tm[536] = 4695;
assign te[536] = 13;
assign s[537] = 6258647;
assign tm[537] = 4693;
assign te[537] = 13;
assign s[538] = 6263337;
assign tm[538] = 4692;
assign te[538] = 13;
assign s[539] = 6268027;
assign tm[539] = 4690;
assign te[539] = 13;
assign s[540] = 6272715;
assign tm[540] = 4689;
assign te[540] = 13;
assign s[541] = 6277402;
assign tm[541] = 4687;
assign te[541] = 13;
assign s[542] = 6282086;
assign tm[542] = 4686;
assign te[542] = 13;
assign s[543] = 6286770;
assign tm[543] = 4684;
assign te[543] = 13;
assign s[544] = 6291451;
assign tm[544] = 4683;
assign te[544] = 13;
assign s[545] = 6296132;
assign tm[545] = 4681;
assign te[545] = 13;
assign s[546] = 6300811;
assign tm[546] = 4680;
assign te[546] = 13;
assign s[547] = 6305488;
assign tm[547] = 4678;
assign te[547] = 13;
assign s[548] = 6310164;
assign tm[548] = 4677;
assign te[548] = 13;
assign s[549] = 6314839;
assign tm[549] = 4675;
assign te[549] = 13;
assign s[550] = 6319511;
assign tm[550] = 4674;
assign te[550] = 13;
assign s[551] = 6324183;
assign tm[551] = 4672;
assign te[551] = 13;
assign s[552] = 6328853;
assign tm[552] = 4671;
assign te[552] = 13;
assign s[553] = 6333522;
assign tm[553] = 4669;
assign te[553] = 13;
assign s[554] = 6338189;
assign tm[554] = 4668;
assign te[554] = 13;
assign s[555] = 6342854;
assign tm[555] = 4667;
assign te[555] = 13;
assign s[556] = 6347518;
assign tm[556] = 4665;
assign te[556] = 13;
assign s[557] = 6352181;
assign tm[557] = 4664;
assign te[557] = 13;
assign s[558] = 6356841;
assign tm[558] = 4662;
assign te[558] = 13;
assign s[559] = 6361501;
assign tm[559] = 4661;
assign te[559] = 13;
assign s[560] = 6366159;
assign tm[560] = 4659;
assign te[560] = 13;
assign s[561] = 6370816;
assign tm[561] = 4658;
assign te[561] = 13;
assign s[562] = 6375472;
assign tm[562] = 4656;
assign te[562] = 13;
assign s[563] = 6380124;
assign tm[563] = 4655;
assign te[563] = 13;
assign s[564] = 6384778;
assign tm[564] = 4653;
assign te[564] = 13;
assign s[565] = 6389429;
assign tm[565] = 4652;
assign te[565] = 13;
assign s[566] = 6394078;
assign tm[566] = 4650;
assign te[566] = 13;
assign s[567] = 6398726;
assign tm[567] = 4649;
assign te[567] = 13;
assign s[568] = 6403372;
assign tm[568] = 4647;
assign te[568] = 13;
assign s[569] = 6408018;
assign tm[569] = 4646;
assign te[569] = 13;
assign s[570] = 6412661;
assign tm[570] = 4644;
assign te[570] = 13;
assign s[571] = 6417303;
assign tm[571] = 4643;
assign te[571] = 13;
assign s[572] = 6421944;
assign tm[572] = 4642;
assign te[572] = 13;
assign s[573] = 6426583;
assign tm[573] = 4640;
assign te[573] = 13;
assign s[574] = 6431220;
assign tm[574] = 4639;
assign te[574] = 13;
assign s[575] = 6435857;
assign tm[575] = 4637;
assign te[575] = 13;
assign s[576] = 6440491;
assign tm[576] = 4636;
assign te[576] = 13;
assign s[577] = 6445125;
assign tm[577] = 4634;
assign te[577] = 13;
assign s[578] = 6449757;
assign tm[578] = 4633;
assign te[578] = 13;
assign s[579] = 6454388;
assign tm[579] = 4631;
assign te[579] = 13;
assign s[580] = 6459016;
assign tm[580] = 4630;
assign te[580] = 13;
assign s[581] = 6463644;
assign tm[581] = 4629;
assign te[581] = 13;
assign s[582] = 6468270;
assign tm[582] = 4627;
assign te[582] = 13;
assign s[583] = 6472895;
assign tm[583] = 4626;
assign te[583] = 13;
assign s[584] = 6477518;
assign tm[584] = 4624;
assign te[584] = 13;
assign s[585] = 6482140;
assign tm[585] = 4623;
assign te[585] = 13;
assign s[586] = 6486760;
assign tm[586] = 4621;
assign te[586] = 13;
assign s[587] = 6491379;
assign tm[587] = 4620;
assign te[587] = 13;
assign s[588] = 6495997;
assign tm[588] = 4618;
assign te[588] = 13;
assign s[589] = 6500613;
assign tm[589] = 4617;
assign te[589] = 13;
assign s[590] = 6505227;
assign tm[590] = 4616;
assign te[590] = 13;
assign s[591] = 6509841;
assign tm[591] = 4614;
assign te[591] = 13;
assign s[592] = 6514453;
assign tm[592] = 4613;
assign te[592] = 13;
assign s[593] = 6519063;
assign tm[593] = 4611;
assign te[593] = 13;
assign s[594] = 6523671;
assign tm[594] = 4610;
assign te[594] = 13;
assign s[595] = 6528279;
assign tm[595] = 4608;
assign te[595] = 13;
assign s[596] = 6532885;
assign tm[596] = 4607;
assign te[596] = 13;
assign s[597] = 6537490;
assign tm[597] = 4606;
assign te[597] = 13;
assign s[598] = 6542094;
assign tm[598] = 4604;
assign te[598] = 13;
assign s[599] = 6546695;
assign tm[599] = 4603;
assign te[599] = 13;
assign s[600] = 6551296;
assign tm[600] = 4601;
assign te[600] = 13;
assign s[601] = 6555895;
assign tm[601] = 4600;
assign te[601] = 13;
assign s[602] = 6560492;
assign tm[602] = 4599;
assign te[602] = 13;
assign s[603] = 6565089;
assign tm[603] = 4597;
assign te[603] = 13;
assign s[604] = 6569683;
assign tm[604] = 4596;
assign te[604] = 13;
assign s[605] = 6574277;
assign tm[605] = 4594;
assign te[605] = 13;
assign s[606] = 6578868;
assign tm[606] = 4593;
assign te[606] = 13;
assign s[607] = 6583459;
assign tm[607] = 4591;
assign te[607] = 13;
assign s[608] = 6588048;
assign tm[608] = 4590;
assign te[608] = 13;
assign s[609] = 6592636;
assign tm[609] = 4589;
assign te[609] = 13;
assign s[610] = 6597222;
assign tm[610] = 4587;
assign te[610] = 13;
assign s[611] = 6601807;
assign tm[611] = 4586;
assign te[611] = 13;
assign s[612] = 6606390;
assign tm[612] = 4584;
assign te[612] = 13;
assign s[613] = 6610973;
assign tm[613] = 4583;
assign te[613] = 13;
assign s[614] = 6615554;
assign tm[614] = 4582;
assign te[614] = 13;
assign s[615] = 6620133;
assign tm[615] = 4580;
assign te[615] = 13;
assign s[616] = 6624711;
assign tm[616] = 4579;
assign te[616] = 13;
assign s[617] = 6629287;
assign tm[617] = 4577;
assign te[617] = 13;
assign s[618] = 6633862;
assign tm[618] = 4576;
assign te[618] = 13;
assign s[619] = 6638437;
assign tm[619] = 4575;
assign te[619] = 13;
assign s[620] = 6643009;
assign tm[620] = 4573;
assign te[620] = 13;
assign s[621] = 6647580;
assign tm[621] = 4572;
assign te[621] = 13;
assign s[622] = 6652150;
assign tm[622] = 4570;
assign te[622] = 13;
assign s[623] = 6656718;
assign tm[623] = 4569;
assign te[623] = 13;
assign s[624] = 6661285;
assign tm[624] = 4568;
assign te[624] = 13;
assign s[625] = 6665850;
assign tm[625] = 4566;
assign te[625] = 13;
assign s[626] = 6670414;
assign tm[626] = 4565;
assign te[626] = 13;
assign s[627] = 6674977;
assign tm[627] = 4564;
assign te[627] = 13;
assign s[628] = 6679538;
assign tm[628] = 4562;
assign te[628] = 13;
assign s[629] = 6684098;
assign tm[629] = 4561;
assign te[629] = 13;
assign s[630] = 6688656;
assign tm[630] = 4559;
assign te[630] = 13;
assign s[631] = 6693214;
assign tm[631] = 4558;
assign te[631] = 13;
assign s[632] = 6697769;
assign tm[632] = 4557;
assign te[632] = 13;
assign s[633] = 6702324;
assign tm[633] = 4555;
assign te[633] = 13;
assign s[634] = 6706877;
assign tm[634] = 4554;
assign te[634] = 13;
assign s[635] = 6711429;
assign tm[635] = 4553;
assign te[635] = 13;
assign s[636] = 6715978;
assign tm[636] = 4551;
assign te[636] = 13;
assign s[637] = 6720527;
assign tm[637] = 4550;
assign te[637] = 13;
assign s[638] = 6725075;
assign tm[638] = 4548;
assign te[638] = 13;
assign s[639] = 6729620;
assign tm[639] = 4547;
assign te[639] = 13;
assign s[640] = 6734166;
assign tm[640] = 4546;
assign te[640] = 13;
assign s[641] = 6738709;
assign tm[641] = 4544;
assign te[641] = 13;
assign s[642] = 6743250;
assign tm[642] = 4543;
assign te[642] = 13;
assign s[643] = 6747792;
assign tm[643] = 4542;
assign te[643] = 13;
assign s[644] = 6752331;
assign tm[644] = 4540;
assign te[644] = 13;
assign s[645] = 6756869;
assign tm[645] = 4539;
assign te[645] = 13;
assign s[646] = 6761405;
assign tm[646] = 4537;
assign te[646] = 13;
assign s[647] = 6765941;
assign tm[647] = 4536;
assign te[647] = 13;
assign s[648] = 6770475;
assign tm[648] = 4535;
assign te[648] = 13;
assign s[649] = 6775008;
assign tm[649] = 4533;
assign te[649] = 13;
assign s[650] = 6779539;
assign tm[650] = 4532;
assign te[650] = 13;
assign s[651] = 6784068;
assign tm[651] = 4531;
assign te[651] = 13;
assign s[652] = 6788597;
assign tm[652] = 4529;
assign te[652] = 13;
assign s[653] = 6793125;
assign tm[653] = 4528;
assign te[653] = 13;
assign s[654] = 6797649;
assign tm[654] = 4527;
assign te[654] = 13;
assign s[655] = 6802174;
assign tm[655] = 4525;
assign te[655] = 13;
assign s[656] = 6806697;
assign tm[656] = 4524;
assign te[656] = 13;
assign s[657] = 6811219;
assign tm[657] = 4523;
assign te[657] = 13;
assign s[658] = 6815739;
assign tm[658] = 4521;
assign te[658] = 13;
assign s[659] = 6820259;
assign tm[659] = 4520;
assign te[659] = 13;
assign s[660] = 6824776;
assign tm[660] = 4519;
assign te[660] = 13;
assign s[661] = 6829292;
assign tm[661] = 4517;
assign te[661] = 13;
assign s[662] = 6833807;
assign tm[662] = 4516;
assign te[662] = 13;
assign s[663] = 6838321;
assign tm[663] = 4515;
assign te[663] = 13;
assign s[664] = 6842834;
assign tm[664] = 4513;
assign te[664] = 13;
assign s[665] = 6847345;
assign tm[665] = 4512;
assign te[665] = 13;
assign s[666] = 6851854;
assign tm[666] = 4511;
assign te[666] = 13;
assign s[667] = 6856363;
assign tm[667] = 4509;
assign te[667] = 13;
assign s[668] = 6860869;
assign tm[668] = 4508;
assign te[668] = 13;
assign s[669] = 6865375;
assign tm[669] = 4507;
assign te[669] = 13;
assign s[670] = 6869880;
assign tm[670] = 4505;
assign te[670] = 13;
assign s[671] = 6874383;
assign tm[671] = 4504;
assign te[671] = 13;
assign s[672] = 6878884;
assign tm[672] = 4503;
assign te[672] = 13;
assign s[673] = 6883385;
assign tm[673] = 4501;
assign te[673] = 13;
assign s[674] = 6887884;
assign tm[674] = 4500;
assign te[674] = 13;
assign s[675] = 6892381;
assign tm[675] = 4499;
assign te[675] = 13;
assign s[676] = 6896878;
assign tm[676] = 4497;
assign te[676] = 13;
assign s[677] = 6901373;
assign tm[677] = 4496;
assign te[677] = 13;
assign s[678] = 6905866;
assign tm[678] = 4495;
assign te[678] = 13;
assign s[679] = 6910359;
assign tm[679] = 4493;
assign te[679] = 13;
assign s[680] = 6914851;
assign tm[680] = 4492;
assign te[680] = 13;
assign s[681] = 6919340;
assign tm[681] = 4491;
assign te[681] = 13;
assign s[682] = 6923828;
assign tm[682] = 4489;
assign te[682] = 13;
assign s[683] = 6928316;
assign tm[683] = 4488;
assign te[683] = 13;
assign s[684] = 6932802;
assign tm[684] = 4487;
assign te[684] = 13;
assign s[685] = 6937286;
assign tm[685] = 4485;
assign te[685] = 13;
assign s[686] = 6941770;
assign tm[686] = 4484;
assign te[686] = 13;
assign s[687] = 6946251;
assign tm[687] = 4483;
assign te[687] = 13;
assign s[688] = 6950732;
assign tm[688] = 4481;
assign te[688] = 13;
assign s[689] = 6955212;
assign tm[689] = 4480;
assign te[689] = 13;
assign s[690] = 6959689;
assign tm[690] = 4479;
assign te[690] = 13;
assign s[691] = 6964166;
assign tm[691] = 4477;
assign te[691] = 13;
assign s[692] = 6968641;
assign tm[692] = 4476;
assign te[692] = 13;
assign s[693] = 6973114;
assign tm[693] = 4475;
assign te[693] = 13;
assign s[694] = 6977588;
assign tm[694] = 4474;
assign te[694] = 13;
assign s[695] = 6982060;
assign tm[695] = 4472;
assign te[695] = 13;
assign s[696] = 6986529;
assign tm[696] = 4471;
assign te[696] = 13;
assign s[697] = 6990999;
assign tm[697] = 4470;
assign te[697] = 13;
assign s[698] = 6995467;
assign tm[698] = 4468;
assign te[698] = 13;
assign s[699] = 6999932;
assign tm[699] = 4467;
assign te[699] = 13;
assign s[700] = 7004398;
assign tm[700] = 4466;
assign te[700] = 13;
assign s[701] = 7008861;
assign tm[701] = 4464;
assign te[701] = 13;
assign s[702] = 7013324;
assign tm[702] = 4463;
assign te[702] = 13;
assign s[703] = 7017785;
assign tm[703] = 4462;
assign te[703] = 13;
assign s[704] = 7022244;
assign tm[704] = 4461;
assign te[704] = 13;
assign s[705] = 7026703;
assign tm[705] = 4459;
assign te[705] = 13;
assign s[706] = 7031160;
assign tm[706] = 4458;
assign te[706] = 13;
assign s[707] = 7035617;
assign tm[707] = 4457;
assign te[707] = 13;
assign s[708] = 7040071;
assign tm[708] = 4455;
assign te[708] = 13;
assign s[709] = 7044524;
assign tm[709] = 4454;
assign te[709] = 13;
assign s[710] = 7048977;
assign tm[710] = 4453;
assign te[710] = 13;
assign s[711] = 7053428;
assign tm[711] = 4452;
assign te[711] = 13;
assign s[712] = 7057876;
assign tm[712] = 4450;
assign te[712] = 13;
assign s[713] = 7062325;
assign tm[713] = 4449;
assign te[713] = 13;
assign s[714] = 7066772;
assign tm[714] = 4448;
assign te[714] = 13;
assign s[715] = 7071217;
assign tm[715] = 4446;
assign te[715] = 13;
assign s[716] = 7075662;
assign tm[716] = 4445;
assign te[716] = 13;
assign s[717] = 7080104;
assign tm[717] = 4444;
assign te[717] = 13;
assign s[718] = 7084547;
assign tm[718] = 4443;
assign te[718] = 13;
assign s[719] = 7088987;
assign tm[719] = 4441;
assign te[719] = 13;
assign s[720] = 7093426;
assign tm[720] = 4440;
assign te[720] = 13;
assign s[721] = 7097865;
assign tm[721] = 4439;
assign te[721] = 13;
assign s[722] = 7102302;
assign tm[722] = 4438;
assign te[722] = 13;
assign s[723] = 7106737;
assign tm[723] = 4436;
assign te[723] = 13;
assign s[724] = 7111171;
assign tm[724] = 4435;
assign te[724] = 13;
assign s[725] = 7115604;
assign tm[725] = 4434;
assign te[725] = 13;
assign s[726] = 7120036;
assign tm[726] = 4432;
assign te[726] = 13;
assign s[727] = 7124466;
assign tm[727] = 4431;
assign te[727] = 13;
assign s[728] = 7128896;
assign tm[728] = 4430;
assign te[728] = 13;
assign s[729] = 7133323;
assign tm[729] = 4429;
assign te[729] = 13;
assign s[730] = 7137750;
assign tm[730] = 4427;
assign te[730] = 13;
assign s[731] = 7142176;
assign tm[731] = 4426;
assign te[731] = 13;
assign s[732] = 7146599;
assign tm[732] = 4425;
assign te[732] = 13;
assign s[733] = 7151022;
assign tm[733] = 4424;
assign te[733] = 13;
assign s[734] = 7155444;
assign tm[734] = 4422;
assign te[734] = 13;
assign s[735] = 7159864;
assign tm[735] = 4421;
assign te[735] = 13;
assign s[736] = 7164284;
assign tm[736] = 4420;
assign te[736] = 13;
assign s[737] = 7168701;
assign tm[737] = 4419;
assign te[737] = 13;
assign s[738] = 7173118;
assign tm[738] = 4417;
assign te[738] = 13;
assign s[739] = 7177532;
assign tm[739] = 4416;
assign te[739] = 13;
assign s[740] = 7181946;
assign tm[740] = 4415;
assign te[740] = 13;
assign s[741] = 7186360;
assign tm[741] = 4414;
assign te[741] = 13;
assign s[742] = 7190772;
assign tm[742] = 4412;
assign te[742] = 13;
assign s[743] = 7195181;
assign tm[743] = 4411;
assign te[743] = 13;
assign s[744] = 7199590;
assign tm[744] = 4410;
assign te[744] = 13;
assign s[745] = 7203998;
assign tm[745] = 4409;
assign te[745] = 13;
assign s[746] = 7208405;
assign tm[746] = 4407;
assign te[746] = 13;
assign s[747] = 7212810;
assign tm[747] = 4406;
assign te[747] = 13;
assign s[748] = 7217214;
assign tm[748] = 4405;
assign te[748] = 13;
assign s[749] = 7221617;
assign tm[749] = 4404;
assign te[749] = 13;
assign s[750] = 7226019;
assign tm[750] = 4402;
assign te[750] = 13;
assign s[751] = 7230419;
assign tm[751] = 4401;
assign te[751] = 13;
assign s[752] = 7234818;
assign tm[752] = 4400;
assign te[752] = 13;
assign s[753] = 7239216;
assign tm[753] = 4399;
assign te[753] = 13;
assign s[754] = 7243613;
assign tm[754] = 4397;
assign te[754] = 13;
assign s[755] = 7248008;
assign tm[755] = 4396;
assign te[755] = 13;
assign s[756] = 7252402;
assign tm[756] = 4395;
assign te[756] = 13;
assign s[757] = 7256795;
assign tm[757] = 4394;
assign te[757] = 13;
assign s[758] = 7261187;
assign tm[758] = 4392;
assign te[758] = 13;
assign s[759] = 7265577;
assign tm[759] = 4391;
assign te[759] = 13;
assign s[760] = 7269967;
assign tm[760] = 4390;
assign te[760] = 13;
assign s[761] = 7274354;
assign tm[761] = 4389;
assign te[761] = 13;
assign s[762] = 7278741;
assign tm[762] = 4387;
assign te[762] = 13;
assign s[763] = 7283127;
assign tm[763] = 4386;
assign te[763] = 13;
assign s[764] = 7287510;
assign tm[764] = 4385;
assign te[764] = 13;
assign s[765] = 7291893;
assign tm[765] = 4384;
assign te[765] = 13;
assign s[766] = 7296276;
assign tm[766] = 4383;
assign te[766] = 13;
assign s[767] = 7300657;
assign tm[767] = 4381;
assign te[767] = 13;
assign s[768] = 7305036;
assign tm[768] = 4380;
assign te[768] = 13;
assign s[769] = 7309414;
assign tm[769] = 4379;
assign te[769] = 13;
assign s[770] = 7313791;
assign tm[770] = 4378;
assign te[770] = 13;
assign s[771] = 7318168;
assign tm[771] = 4376;
assign te[771] = 13;
assign s[772] = 7322542;
assign tm[772] = 4375;
assign te[772] = 13;
assign s[773] = 7326915;
assign tm[773] = 4374;
assign te[773] = 13;
assign s[774] = 7331287;
assign tm[774] = 4373;
assign te[774] = 13;
assign s[775] = 7335657;
assign tm[775] = 4372;
assign te[775] = 13;
assign s[776] = 7340028;
assign tm[776] = 4370;
assign te[776] = 13;
assign s[777] = 7344397;
assign tm[777] = 4369;
assign te[777] = 13;
assign s[778] = 7348763;
assign tm[778] = 4368;
assign te[778] = 13;
assign s[779] = 7353130;
assign tm[779] = 4367;
assign te[779] = 13;
assign s[780] = 7357494;
assign tm[780] = 4366;
assign te[780] = 13;
assign s[781] = 7361857;
assign tm[781] = 4364;
assign te[781] = 13;
assign s[782] = 7366220;
assign tm[782] = 4363;
assign te[782] = 13;
assign s[783] = 7370582;
assign tm[783] = 4362;
assign te[783] = 13;
assign s[784] = 7374941;
assign tm[784] = 4361;
assign te[784] = 13;
assign s[785] = 7379300;
assign tm[785] = 4359;
assign te[785] = 13;
assign s[786] = 7383657;
assign tm[786] = 4358;
assign te[786] = 13;
assign s[787] = 7388014;
assign tm[787] = 4357;
assign te[787] = 13;
assign s[788] = 7392369;
assign tm[788] = 4356;
assign te[788] = 13;
assign s[789] = 7396723;
assign tm[789] = 4355;
assign te[789] = 13;
assign s[790] = 7401077;
assign tm[790] = 4353;
assign te[790] = 13;
assign s[791] = 7405428;
assign tm[791] = 4352;
assign te[791] = 13;
assign s[792] = 7409777;
assign tm[792] = 4351;
assign te[792] = 13;
assign s[793] = 7414127;
assign tm[793] = 4350;
assign te[793] = 13;
assign s[794] = 7418476;
assign tm[794] = 4349;
assign te[794] = 13;
assign s[795] = 7422822;
assign tm[795] = 4347;
assign te[795] = 13;
assign s[796] = 7427168;
assign tm[796] = 4346;
assign te[796] = 13;
assign s[797] = 7431512;
assign tm[797] = 4345;
assign te[797] = 13;
assign s[798] = 7435856;
assign tm[798] = 4344;
assign te[798] = 13;
assign s[799] = 7440198;
assign tm[799] = 4343;
assign te[799] = 13;
assign s[800] = 7444538;
assign tm[800] = 4342;
assign te[800] = 13;
assign s[801] = 7448877;
assign tm[801] = 4340;
assign te[801] = 13;
assign s[802] = 7453216;
assign tm[802] = 4339;
assign te[802] = 13;
assign s[803] = 7457553;
assign tm[803] = 4338;
assign te[803] = 13;
assign s[804] = 7461889;
assign tm[804] = 4337;
assign te[804] = 13;
assign s[805] = 7466224;
assign tm[805] = 4336;
assign te[805] = 13;
assign s[806] = 7470557;
assign tm[806] = 4334;
assign te[806] = 13;
assign s[807] = 7474890;
assign tm[807] = 4333;
assign te[807] = 13;
assign s[808] = 7479222;
assign tm[808] = 4332;
assign te[808] = 13;
assign s[809] = 7483552;
assign tm[809] = 4331;
assign te[809] = 13;
assign s[810] = 7487881;
assign tm[810] = 4330;
assign te[810] = 13;
assign s[811] = 7492209;
assign tm[811] = 4328;
assign te[811] = 13;
assign s[812] = 7496535;
assign tm[812] = 4327;
assign te[812] = 13;
assign s[813] = 7500860;
assign tm[813] = 4326;
assign te[813] = 13;
assign s[814] = 7505185;
assign tm[814] = 4325;
assign te[814] = 13;
assign s[815] = 7509508;
assign tm[815] = 4324;
assign te[815] = 13;
assign s[816] = 7513830;
assign tm[816] = 4323;
assign te[816] = 13;
assign s[817] = 7518150;
assign tm[817] = 4321;
assign te[817] = 13;
assign s[818] = 7522471;
assign tm[818] = 4320;
assign te[818] = 13;
assign s[819] = 7526789;
assign tm[819] = 4319;
assign te[819] = 13;
assign s[820] = 7531106;
assign tm[820] = 4318;
assign te[820] = 13;
assign s[821] = 7535422;
assign tm[821] = 4317;
assign te[821] = 13;
assign s[822] = 7539737;
assign tm[822] = 4316;
assign te[822] = 13;
assign s[823] = 7544050;
assign tm[823] = 4314;
assign te[823] = 13;
assign s[824] = 7548363;
assign tm[824] = 4313;
assign te[824] = 13;
assign s[825] = 7552674;
assign tm[825] = 4312;
assign te[825] = 13;
assign s[826] = 7556984;
assign tm[826] = 4311;
assign te[826] = 13;
assign s[827] = 7561294;
assign tm[827] = 4310;
assign te[827] = 13;
assign s[828] = 7565601;
assign tm[828] = 4309;
assign te[828] = 13;
assign s[829] = 7569908;
assign tm[829] = 4307;
assign te[829] = 13;
assign s[830] = 7574214;
assign tm[830] = 4306;
assign te[830] = 13;
assign s[831] = 7578518;
assign tm[831] = 4305;
assign te[831] = 13;
assign s[832] = 7582822;
assign tm[832] = 4304;
assign te[832] = 13;
assign s[833] = 7587124;
assign tm[833] = 4303;
assign te[833] = 13;
assign s[834] = 7591424;
assign tm[834] = 4302;
assign te[834] = 13;
assign s[835] = 7595724;
assign tm[835] = 4300;
assign te[835] = 13;
assign s[836] = 7600022;
assign tm[836] = 4299;
assign te[836] = 13;
assign s[837] = 7604320;
assign tm[837] = 4298;
assign te[837] = 13;
assign s[838] = 7608616;
assign tm[838] = 4297;
assign te[838] = 13;
assign s[839] = 7612913;
assign tm[839] = 4296;
assign te[839] = 13;
assign s[840] = 7617206;
assign tm[840] = 4295;
assign te[840] = 13;
assign s[841] = 7621499;
assign tm[841] = 4293;
assign te[841] = 13;
assign s[842] = 7625790;
assign tm[842] = 4292;
assign te[842] = 13;
assign s[843] = 7630080;
assign tm[843] = 4291;
assign te[843] = 13;
assign s[844] = 7634370;
assign tm[844] = 4290;
assign te[844] = 13;
assign s[845] = 7638658;
assign tm[845] = 4289;
assign te[845] = 13;
assign s[846] = 7642945;
assign tm[846] = 4288;
assign te[846] = 13;
assign s[847] = 7647231;
assign tm[847] = 4287;
assign te[847] = 13;
assign s[848] = 7651517;
assign tm[848] = 4285;
assign te[848] = 13;
assign s[849] = 7655799;
assign tm[849] = 4284;
assign te[849] = 13;
assign s[850] = 7660082;
assign tm[850] = 4283;
assign te[850] = 13;
assign s[851] = 7664364;
assign tm[851] = 4282;
assign te[851] = 13;
assign s[852] = 7668643;
assign tm[852] = 4281;
assign te[852] = 13;
assign s[853] = 7672923;
assign tm[853] = 4280;
assign te[853] = 13;
assign s[854] = 7677201;
assign tm[854] = 4279;
assign te[854] = 13;
assign s[855] = 7681478;
assign tm[855] = 4277;
assign te[855] = 13;
assign s[856] = 7685753;
assign tm[856] = 4276;
assign te[856] = 13;
assign s[857] = 7690027;
assign tm[857] = 4275;
assign te[857] = 13;
assign s[858] = 7694302;
assign tm[858] = 4274;
assign te[858] = 13;
assign s[859] = 7698573;
assign tm[859] = 4273;
assign te[859] = 13;
assign s[860] = 7702846;
assign tm[860] = 4272;
assign te[860] = 13;
assign s[861] = 7707115;
assign tm[861] = 4271;
assign te[861] = 13;
assign s[862] = 7711384;
assign tm[862] = 4269;
assign te[862] = 13;
assign s[863] = 7715652;
assign tm[863] = 4268;
assign te[863] = 13;
assign s[864] = 7719918;
assign tm[864] = 4267;
assign te[864] = 13;
assign s[865] = 7724184;
assign tm[865] = 4266;
assign te[865] = 13;
assign s[866] = 7728448;
assign tm[866] = 4265;
assign te[866] = 13;
assign s[867] = 7732711;
assign tm[867] = 4264;
assign te[867] = 13;
assign s[868] = 7736974;
assign tm[868] = 4263;
assign te[868] = 13;
assign s[869] = 7741235;
assign tm[869] = 4262;
assign te[869] = 13;
assign s[870] = 7745494;
assign tm[870] = 4260;
assign te[870] = 13;
assign s[871] = 7749752;
assign tm[871] = 4259;
assign te[871] = 13;
assign s[872] = 7754009;
assign tm[872] = 4258;
assign te[872] = 13;
assign s[873] = 7758266;
assign tm[873] = 4257;
assign te[873] = 13;
assign s[874] = 7762522;
assign tm[874] = 4256;
assign te[874] = 13;
assign s[875] = 7766775;
assign tm[875] = 4255;
assign te[875] = 13;
assign s[876] = 7771029;
assign tm[876] = 4254;
assign te[876] = 13;
assign s[877] = 7775281;
assign tm[877] = 4253;
assign te[877] = 13;
assign s[878] = 7779532;
assign tm[878] = 4251;
assign te[878] = 13;
assign s[879] = 7783782;
assign tm[879] = 4250;
assign te[879] = 13;
assign s[880] = 7788030;
assign tm[880] = 4249;
assign te[880] = 13;
assign s[881] = 7792278;
assign tm[881] = 4248;
assign te[881] = 13;
assign s[882] = 7796524;
assign tm[882] = 4247;
assign te[882] = 13;
assign s[883] = 7800770;
assign tm[883] = 4246;
assign te[883] = 13;
assign s[884] = 7805014;
assign tm[884] = 4245;
assign te[884] = 13;
assign s[885] = 7809257;
assign tm[885] = 4244;
assign te[885] = 13;
assign s[886] = 7813498;
assign tm[886] = 4243;
assign te[886] = 13;
assign s[887] = 7817739;
assign tm[887] = 4241;
assign te[887] = 13;
assign s[888] = 7821979;
assign tm[888] = 4240;
assign te[888] = 13;
assign s[889] = 7826217;
assign tm[889] = 4239;
assign te[889] = 13;
assign s[890] = 7830456;
assign tm[890] = 4238;
assign te[890] = 13;
assign s[891] = 7834691;
assign tm[891] = 4237;
assign te[891] = 13;
assign s[892] = 7838928;
assign tm[892] = 4236;
assign te[892] = 13;
assign s[893] = 7843163;
assign tm[893] = 4235;
assign te[893] = 13;
assign s[894] = 7847394;
assign tm[894] = 4234;
assign te[894] = 13;
assign s[895] = 7851626;
assign tm[895] = 4233;
assign te[895] = 13;
assign s[896] = 7855858;
assign tm[896] = 4231;
assign te[896] = 13;
assign s[897] = 7860087;
assign tm[897] = 4230;
assign te[897] = 13;
assign s[898] = 7864316;
assign tm[898] = 4229;
assign te[898] = 13;
assign s[899] = 7868543;
assign tm[899] = 4228;
assign te[899] = 13;
assign s[900] = 7872769;
assign tm[900] = 4227;
assign te[900] = 13;
assign s[901] = 7876995;
assign tm[901] = 4226;
assign te[901] = 13;
assign s[902] = 7881219;
assign tm[902] = 4225;
assign te[902] = 13;
assign s[903] = 7885442;
assign tm[903] = 4224;
assign te[903] = 13;
assign s[904] = 7889664;
assign tm[904] = 4223;
assign te[904] = 13;
assign s[905] = 7893886;
assign tm[905] = 4222;
assign te[905] = 13;
assign s[906] = 7898105;
assign tm[906] = 4220;
assign te[906] = 13;
assign s[907] = 7902324;
assign tm[907] = 4219;
assign te[907] = 13;
assign s[908] = 7906543;
assign tm[908] = 4218;
assign te[908] = 13;
assign s[909] = 7910759;
assign tm[909] = 4217;
assign te[909] = 13;
assign s[910] = 7914974;
assign tm[910] = 4216;
assign te[910] = 13;
assign s[911] = 7919189;
assign tm[911] = 4215;
assign te[911] = 13;
assign s[912] = 7923403;
assign tm[912] = 4214;
assign te[912] = 13;
assign s[913] = 7927614;
assign tm[913] = 4213;
assign te[913] = 13;
assign s[914] = 7931825;
assign tm[914] = 4212;
assign te[914] = 13;
assign s[915] = 7936035;
assign tm[915] = 4211;
assign te[915] = 13;
assign s[916] = 7940244;
assign tm[916] = 4210;
assign te[916] = 13;
assign s[917] = 7944453;
assign tm[917] = 4209;
assign te[917] = 13;
assign s[918] = 7948659;
assign tm[918] = 4207;
assign te[918] = 13;
assign s[919] = 7952866;
assign tm[919] = 4206;
assign te[919] = 13;
assign s[920] = 7957070;
assign tm[920] = 4205;
assign te[920] = 13;
assign s[921] = 7961274;
assign tm[921] = 4204;
assign te[921] = 13;
assign s[922] = 7965476;
assign tm[922] = 4203;
assign te[922] = 13;
assign s[923] = 7969678;
assign tm[923] = 4202;
assign te[923] = 13;
assign s[924] = 7973877;
assign tm[924] = 4201;
assign te[924] = 13;
assign s[925] = 7978077;
assign tm[925] = 4200;
assign te[925] = 13;
assign s[926] = 7982275;
assign tm[926] = 4199;
assign te[926] = 13;
assign s[927] = 7986472;
assign tm[927] = 4198;
assign te[927] = 13;
assign s[928] = 7990669;
assign tm[928] = 4197;
assign te[928] = 13;
assign s[929] = 7994864;
assign tm[929] = 4196;
assign te[929] = 13;
assign s[930] = 7999056;
assign tm[930] = 4194;
assign te[930] = 13;
assign s[931] = 8003249;
assign tm[931] = 4193;
assign te[931] = 13;
assign s[932] = 8007442;
assign tm[932] = 4192;
assign te[932] = 13;
assign s[933] = 8011632;
assign tm[933] = 4191;
assign te[933] = 13;
assign s[934] = 8015823;
assign tm[934] = 4190;
assign te[934] = 13;
assign s[935] = 8020010;
assign tm[935] = 4189;
assign te[935] = 13;
assign s[936] = 8024197;
assign tm[936] = 4188;
assign te[936] = 13;
assign s[937] = 8028384;
assign tm[937] = 4187;
assign te[937] = 13;
assign s[938] = 8032570;
assign tm[938] = 4186;
assign te[938] = 13;
assign s[939] = 8036754;
assign tm[939] = 4185;
assign te[939] = 13;
assign s[940] = 8040937;
assign tm[940] = 4184;
assign te[940] = 13;
assign s[941] = 8045120;
assign tm[941] = 4183;
assign te[941] = 13;
assign s[942] = 8049301;
assign tm[942] = 4182;
assign te[942] = 13;
assign s[943] = 8053480;
assign tm[943] = 4181;
assign te[943] = 13;
assign s[944] = 8057660;
assign tm[944] = 4180;
assign te[944] = 13;
assign s[945] = 8061837;
assign tm[945] = 4178;
assign te[945] = 13;
assign s[946] = 8066014;
assign tm[946] = 4177;
assign te[946] = 13;
assign s[947] = 8070190;
assign tm[947] = 4176;
assign te[947] = 13;
assign s[948] = 8074365;
assign tm[948] = 4175;
assign te[948] = 13;
assign s[949] = 8078538;
assign tm[949] = 4174;
assign te[949] = 13;
assign s[950] = 8082711;
assign tm[950] = 4173;
assign te[950] = 13;
assign s[951] = 8086882;
assign tm[951] = 4172;
assign te[951] = 13;
assign s[952] = 8091054;
assign tm[952] = 4171;
assign te[952] = 13;
assign s[953] = 8095223;
assign tm[953] = 4170;
assign te[953] = 13;
assign s[954] = 8099391;
assign tm[954] = 4169;
assign te[954] = 13;
assign s[955] = 8103558;
assign tm[955] = 4168;
assign te[955] = 13;
assign s[956] = 8107725;
assign tm[956] = 4167;
assign te[956] = 13;
assign s[957] = 8111889;
assign tm[957] = 4166;
assign te[957] = 13;
assign s[958] = 8116054;
assign tm[958] = 4165;
assign te[958] = 13;
assign s[959] = 8120216;
assign tm[959] = 4164;
assign te[959] = 13;
assign s[960] = 8124378;
assign tm[960] = 4163;
assign te[960] = 13;
assign s[961] = 8128540;
assign tm[961] = 4162;
assign te[961] = 13;
assign s[962] = 8132700;
assign tm[962] = 4161;
assign te[962] = 13;
assign s[963] = 8136859;
assign tm[963] = 4159;
assign te[963] = 13;
assign s[964] = 8141017;
assign tm[964] = 4158;
assign te[964] = 13;
assign s[965] = 8145174;
assign tm[965] = 4157;
assign te[965] = 13;
assign s[966] = 8149330;
assign tm[966] = 4156;
assign te[966] = 13;
assign s[967] = 8153485;
assign tm[967] = 4155;
assign te[967] = 13;
assign s[968] = 8157638;
assign tm[968] = 4154;
assign te[968] = 13;
assign s[969] = 8161790;
assign tm[969] = 4153;
assign te[969] = 13;
assign s[970] = 8165942;
assign tm[970] = 4152;
assign te[970] = 13;
assign s[971] = 8170093;
assign tm[971] = 4151;
assign te[971] = 13;
assign s[972] = 8174242;
assign tm[972] = 4150;
assign te[972] = 13;
assign s[973] = 8178391;
assign tm[973] = 4149;
assign te[973] = 13;
assign s[974] = 8182539;
assign tm[974] = 4148;
assign te[974] = 13;
assign s[975] = 8186685;
assign tm[975] = 4147;
assign te[975] = 13;
assign s[976] = 8190830;
assign tm[976] = 4146;
assign te[976] = 13;
assign s[977] = 8194975;
assign tm[977] = 4145;
assign te[977] = 13;
assign s[978] = 8199117;
assign tm[978] = 4144;
assign te[978] = 13;
assign s[979] = 8203260;
assign tm[979] = 4143;
assign te[979] = 13;
assign s[980] = 8207400;
assign tm[980] = 4142;
assign te[980] = 13;
assign s[981] = 8211541;
assign tm[981] = 4141;
assign te[981] = 13;
assign s[982] = 8215681;
assign tm[982] = 4140;
assign te[982] = 13;
assign s[983] = 8219819;
assign tm[983] = 4139;
assign te[983] = 13;
assign s[984] = 8223956;
assign tm[984] = 4138;
assign te[984] = 13;
assign s[985] = 8228092;
assign tm[985] = 4137;
assign te[985] = 13;
assign s[986] = 8232227;
assign tm[986] = 4136;
assign te[986] = 13;
assign s[987] = 8236362;
assign tm[987] = 4135;
assign te[987] = 13;
assign s[988] = 8240494;
assign tm[988] = 4134;
assign te[988] = 13;
assign s[989] = 8244626;
assign tm[989] = 4132;
assign te[989] = 13;
assign s[990] = 8248757;
assign tm[990] = 4131;
assign te[990] = 13;
assign s[991] = 8252887;
assign tm[991] = 4130;
assign te[991] = 13;
assign s[992] = 8257015;
assign tm[992] = 4129;
assign te[992] = 13;
assign s[993] = 8261143;
assign tm[993] = 4128;
assign te[993] = 13;
assign s[994] = 8265270;
assign tm[994] = 4127;
assign te[994] = 13;
assign s[995] = 8269396;
assign tm[995] = 4126;
assign te[995] = 13;
assign s[996] = 8273521;
assign tm[996] = 4125;
assign te[996] = 13;
assign s[997] = 8277645;
assign tm[997] = 4124;
assign te[997] = 13;
assign s[998] = 8281767;
assign tm[998] = 4123;
assign te[998] = 13;
assign s[999] = 8285888;
assign tm[999] = 4122;
assign te[999] = 13;
assign s[1000] = 8290010;
assign tm[1000] = 4121;
assign te[1000] = 13;
assign s[1001] = 8294130;
assign tm[1001] = 4120;
assign te[1001] = 13;
assign s[1002] = 8298248;
assign tm[1002] = 4119;
assign te[1002] = 13;
assign s[1003] = 8302366;
assign tm[1003] = 4118;
assign te[1003] = 13;
assign s[1004] = 8306482;
assign tm[1004] = 4117;
assign te[1004] = 13;
assign s[1005] = 8310599;
assign tm[1005] = 4116;
assign te[1005] = 13;
assign s[1006] = 8314713;
assign tm[1006] = 4115;
assign te[1006] = 13;
assign s[1007] = 8318826;
assign tm[1007] = 4114;
assign te[1007] = 13;
assign s[1008] = 8322940;
assign tm[1008] = 4113;
assign te[1008] = 13;
assign s[1009] = 8327051;
assign tm[1009] = 4112;
assign te[1009] = 13;
assign s[1010] = 8331162;
assign tm[1010] = 4111;
assign te[1010] = 13;
assign s[1011] = 8335270;
assign tm[1011] = 4110;
assign te[1011] = 13;
assign s[1012] = 8339379;
assign tm[1012] = 4109;
assign te[1012] = 13;
assign s[1013] = 8343487;
assign tm[1013] = 4108;
assign te[1013] = 13;
assign s[1014] = 8347595;
assign tm[1014] = 4107;
assign te[1014] = 13;
assign s[1015] = 8351699;
assign tm[1015] = 4106;
assign te[1015] = 13;
assign s[1016] = 8355804;
assign tm[1016] = 4105;
assign te[1016] = 13;
assign s[1017] = 8359908;
assign tm[1017] = 4104;
assign te[1017] = 13;
assign s[1018] = 8364010;
assign tm[1018] = 4103;
assign te[1018] = 13;
assign s[1019] = 8368112;
assign tm[1019] = 4102;
assign te[1019] = 13;
assign s[1020] = 8372212;
assign tm[1020] = 4101;
assign te[1020] = 13;
assign s[1021] = 8376312;
assign tm[1021] = 4100;
assign te[1021] = 13;
assign s[1022] = 8380410;
assign tm[1022] = 4099;
assign te[1022] = 13;
assign s[1023] = 8384508;
assign tm[1023] = 4098;
assign te[1023] = 13;
assign s[1024] = 0;
assign tm[1024] = 4098;
assign te[1024] = 13;
assign s[1025] = 4090;
assign tm[1025] = 4096;
assign te[1025] = 13;
assign s[1026] = 8183;
assign tm[1026] = 8189;
assign te[1026] = 14;
assign s[1027] = 12274;
assign tm[1027] = 8185;
assign te[1027] = 14;
assign s[1028] = 16364;
assign tm[1028] = 8182;
assign te[1028] = 14;
assign s[1029] = 20450;
assign tm[1029] = 8178;
assign te[1029] = 14;
assign s[1030] = 24536;
assign tm[1030] = 8174;
assign te[1030] = 14;
assign s[1031] = 28618;
assign tm[1031] = 8170;
assign te[1031] = 14;
assign s[1032] = 32699;
assign tm[1032] = 8166;
assign te[1032] = 14;
assign s[1033] = 36779;
assign tm[1033] = 8162;
assign te[1033] = 14;
assign s[1034] = 40856;
assign tm[1034] = 8158;
assign te[1034] = 14;
assign s[1035] = 44931;
assign tm[1035] = 8154;
assign te[1035] = 14;
assign s[1036] = 49004;
assign tm[1036] = 8150;
assign te[1036] = 14;
assign s[1037] = 53075;
assign tm[1037] = 8146;
assign te[1037] = 14;
assign s[1038] = 57145;
assign tm[1038] = 8142;
assign te[1038] = 14;
assign s[1039] = 61212;
assign tm[1039] = 8138;
assign te[1039] = 14;
assign s[1040] = 65277;
assign tm[1040] = 8134;
assign te[1040] = 14;
assign s[1041] = 69341;
assign tm[1041] = 8130;
assign te[1041] = 14;
assign s[1042] = 73402;
assign tm[1042] = 8126;
assign te[1042] = 14;
assign s[1043] = 77462;
assign tm[1043] = 8122;
assign te[1043] = 14;
assign s[1044] = 81519;
assign tm[1044] = 8118;
assign te[1044] = 14;
assign s[1045] = 85574;
assign tm[1045] = 8115;
assign te[1045] = 14;
assign s[1046] = 89628;
assign tm[1046] = 8111;
assign te[1046] = 14;
assign s[1047] = 93680;
assign tm[1047] = 8107;
assign te[1047] = 14;
assign s[1048] = 97730;
assign tm[1048] = 8103;
assign te[1048] = 14;
assign s[1049] = 101777;
assign tm[1049] = 8099;
assign te[1049] = 14;
assign s[1050] = 105824;
assign tm[1050] = 8095;
assign te[1050] = 14;
assign s[1051] = 109868;
assign tm[1051] = 8091;
assign te[1051] = 14;
assign s[1052] = 113910;
assign tm[1052] = 8088;
assign te[1052] = 14;
assign s[1053] = 117950;
assign tm[1053] = 8084;
assign te[1053] = 14;
assign s[1054] = 121988;
assign tm[1054] = 8080;
assign te[1054] = 14;
assign s[1055] = 126025;
assign tm[1055] = 8076;
assign te[1055] = 14;
assign s[1056] = 130059;
assign tm[1056] = 8072;
assign te[1056] = 14;
assign s[1057] = 134092;
assign tm[1057] = 8068;
assign te[1057] = 14;
assign s[1058] = 138122;
assign tm[1058] = 8065;
assign te[1058] = 14;
assign s[1059] = 142151;
assign tm[1059] = 8061;
assign te[1059] = 14;
assign s[1060] = 146177;
assign tm[1060] = 8057;
assign te[1060] = 14;
assign s[1061] = 150202;
assign tm[1061] = 8053;
assign te[1061] = 14;
assign s[1062] = 154226;
assign tm[1062] = 8049;
assign te[1062] = 14;
assign s[1063] = 158247;
assign tm[1063] = 8045;
assign te[1063] = 14;
assign s[1064] = 162266;
assign tm[1064] = 8042;
assign te[1064] = 14;
assign s[1065] = 166283;
assign tm[1065] = 8038;
assign te[1065] = 14;
assign s[1066] = 170298;
assign tm[1066] = 8034;
assign te[1066] = 14;
assign s[1067] = 174312;
assign tm[1067] = 8030;
assign te[1067] = 14;
assign s[1068] = 178324;
assign tm[1068] = 8027;
assign te[1068] = 14;
assign s[1069] = 182334;
assign tm[1069] = 8023;
assign te[1069] = 14;
assign s[1070] = 186341;
assign tm[1070] = 8019;
assign te[1070] = 14;
assign s[1071] = 190347;
assign tm[1071] = 8015;
assign te[1071] = 14;
assign s[1072] = 194352;
assign tm[1072] = 8012;
assign te[1072] = 14;
assign s[1073] = 198354;
assign tm[1073] = 8008;
assign te[1073] = 14;
assign s[1074] = 202355;
assign tm[1074] = 8004;
assign te[1074] = 14;
assign s[1075] = 206353;
assign tm[1075] = 8000;
assign te[1075] = 14;
assign s[1076] = 210350;
assign tm[1076] = 7997;
assign te[1076] = 14;
assign s[1077] = 214345;
assign tm[1077] = 7993;
assign te[1077] = 14;
assign s[1078] = 218337;
assign tm[1078] = 7989;
assign te[1078] = 14;
assign s[1079] = 222329;
assign tm[1079] = 7986;
assign te[1079] = 14;
assign s[1080] = 226318;
assign tm[1080] = 7982;
assign te[1080] = 14;
assign s[1081] = 230306;
assign tm[1081] = 7978;
assign te[1081] = 14;
assign s[1082] = 234291;
assign tm[1082] = 7974;
assign te[1082] = 14;
assign s[1083] = 238275;
assign tm[1083] = 7971;
assign te[1083] = 14;
assign s[1084] = 242257;
assign tm[1084] = 7967;
assign te[1084] = 14;
assign s[1085] = 246237;
assign tm[1085] = 7963;
assign te[1085] = 14;
assign s[1086] = 250215;
assign tm[1086] = 7960;
assign te[1086] = 14;
assign s[1087] = 254192;
assign tm[1087] = 7956;
assign te[1087] = 14;
assign s[1088] = 258167;
assign tm[1088] = 7952;
assign te[1088] = 14;
assign s[1089] = 262140;
assign tm[1089] = 7949;
assign te[1089] = 14;
assign s[1090] = 266110;
assign tm[1090] = 7945;
assign te[1090] = 14;
assign s[1091] = 270079;
assign tm[1091] = 7941;
assign te[1091] = 14;
assign s[1092] = 274047;
assign tm[1092] = 7938;
assign te[1092] = 14;
assign s[1093] = 278012;
assign tm[1093] = 7934;
assign te[1093] = 14;
assign s[1094] = 281976;
assign tm[1094] = 7931;
assign te[1094] = 14;
assign s[1095] = 285938;
assign tm[1095] = 7927;
assign te[1095] = 14;
assign s[1096] = 289898;
assign tm[1096] = 7923;
assign te[1096] = 14;
assign s[1097] = 293856;
assign tm[1097] = 7920;
assign te[1097] = 14;
assign s[1098] = 297813;
assign tm[1098] = 7916;
assign te[1098] = 14;
assign s[1099] = 301767;
assign tm[1099] = 7912;
assign te[1099] = 14;
assign s[1100] = 305721;
assign tm[1100] = 7909;
assign te[1100] = 14;
assign s[1101] = 309671;
assign tm[1101] = 7905;
assign te[1101] = 14;
assign s[1102] = 313621;
assign tm[1102] = 7902;
assign te[1102] = 14;
assign s[1103] = 317568;
assign tm[1103] = 7898;
assign te[1103] = 14;
assign s[1104] = 321514;
assign tm[1104] = 7894;
assign te[1104] = 14;
assign s[1105] = 325458;
assign tm[1105] = 7891;
assign te[1105] = 14;
assign s[1106] = 329400;
assign tm[1106] = 7887;
assign te[1106] = 14;
assign s[1107] = 333340;
assign tm[1107] = 7884;
assign te[1107] = 14;
assign s[1108] = 337279;
assign tm[1108] = 7880;
assign te[1108] = 14;
assign s[1109] = 341216;
assign tm[1109] = 7877;
assign te[1109] = 14;
assign s[1110] = 345151;
assign tm[1110] = 7873;
assign te[1110] = 14;
assign s[1111] = 349084;
assign tm[1111] = 7870;
assign te[1111] = 14;
assign s[1112] = 353015;
assign tm[1112] = 7866;
assign te[1112] = 14;
assign s[1113] = 356945;
assign tm[1113] = 7862;
assign te[1113] = 14;
assign s[1114] = 360873;
assign tm[1114] = 7859;
assign te[1114] = 14;
assign s[1115] = 364799;
assign tm[1115] = 7855;
assign te[1115] = 14;
assign s[1116] = 368723;
assign tm[1116] = 7852;
assign te[1116] = 14;
assign s[1117] = 372646;
assign tm[1117] = 7848;
assign te[1117] = 14;
assign s[1118] = 376567;
assign tm[1118] = 7845;
assign te[1118] = 14;
assign s[1119] = 380487;
assign tm[1119] = 7841;
assign te[1119] = 14;
assign s[1120] = 384403;
assign tm[1120] = 7838;
assign te[1120] = 14;
assign s[1121] = 388319;
assign tm[1121] = 7834;
assign te[1121] = 14;
assign s[1122] = 392233;
assign tm[1122] = 7831;
assign te[1122] = 14;
assign s[1123] = 396145;
assign tm[1123] = 7827;
assign te[1123] = 14;
assign s[1124] = 400056;
assign tm[1124] = 7824;
assign te[1124] = 14;
assign s[1125] = 403964;
assign tm[1125] = 7820;
assign te[1125] = 14;
assign s[1126] = 407871;
assign tm[1126] = 7817;
assign te[1126] = 14;
assign s[1127] = 411777;
assign tm[1127] = 7813;
assign te[1127] = 14;
assign s[1128] = 415680;
assign tm[1128] = 7810;
assign te[1128] = 14;
assign s[1129] = 419581;
assign tm[1129] = 7806;
assign te[1129] = 14;
assign s[1130] = 423482;
assign tm[1130] = 7803;
assign te[1130] = 14;
assign s[1131] = 427380;
assign tm[1131] = 7800;
assign te[1131] = 14;
assign s[1132] = 431277;
assign tm[1132] = 7796;
assign te[1132] = 14;
assign s[1133] = 435172;
assign tm[1133] = 7793;
assign te[1133] = 14;
assign s[1134] = 439065;
assign tm[1134] = 7789;
assign te[1134] = 14;
assign s[1135] = 442956;
assign tm[1135] = 7786;
assign te[1135] = 14;
assign s[1136] = 446846;
assign tm[1136] = 7782;
assign te[1136] = 14;
assign s[1137] = 450734;
assign tm[1137] = 7779;
assign te[1137] = 14;
assign s[1138] = 454620;
assign tm[1138] = 7775;
assign te[1138] = 14;
assign s[1139] = 458504;
assign tm[1139] = 7772;
assign te[1139] = 14;
assign s[1140] = 462388;
assign tm[1140] = 7769;
assign te[1140] = 14;
assign s[1141] = 466269;
assign tm[1141] = 7765;
assign te[1141] = 14;
assign s[1142] = 470148;
assign tm[1142] = 7762;
assign te[1142] = 14;
assign s[1143] = 474026;
assign tm[1143] = 7758;
assign te[1143] = 14;
assign s[1144] = 477902;
assign tm[1144] = 7755;
assign te[1144] = 14;
assign s[1145] = 481776;
assign tm[1145] = 7752;
assign te[1145] = 14;
assign s[1146] = 485649;
assign tm[1146] = 7748;
assign te[1146] = 14;
assign s[1147] = 489520;
assign tm[1147] = 7745;
assign te[1147] = 14;
assign s[1148] = 493389;
assign tm[1148] = 7741;
assign te[1148] = 14;
assign s[1149] = 497257;
assign tm[1149] = 7738;
assign te[1149] = 14;
assign s[1150] = 501123;
assign tm[1150] = 7735;
assign te[1150] = 14;
assign s[1151] = 504987;
assign tm[1151] = 7731;
assign te[1151] = 14;
assign s[1152] = 508850;
assign tm[1152] = 7728;
assign te[1152] = 14;
assign s[1153] = 512711;
assign tm[1153] = 7725;
assign te[1153] = 14;
assign s[1154] = 516570;
assign tm[1154] = 7721;
assign te[1154] = 14;
assign s[1155] = 520428;
assign tm[1155] = 7718;
assign te[1155] = 14;
assign s[1156] = 524283;
assign tm[1156] = 7715;
assign te[1156] = 14;
assign s[1157] = 528137;
assign tm[1157] = 7711;
assign te[1157] = 14;
assign s[1158] = 531991;
assign tm[1158] = 7708;
assign te[1158] = 14;
assign s[1159] = 535841;
assign tm[1159] = 7705;
assign te[1159] = 14;
assign s[1160] = 539690;
assign tm[1160] = 7701;
assign te[1160] = 14;
assign s[1161] = 543538;
assign tm[1161] = 7698;
assign te[1161] = 14;
assign s[1162] = 547384;
assign tm[1162] = 7695;
assign te[1162] = 14;
assign s[1163] = 551228;
assign tm[1163] = 7691;
assign te[1163] = 14;
assign s[1164] = 555071;
assign tm[1164] = 7688;
assign te[1164] = 14;
assign s[1165] = 558911;
assign tm[1165] = 7685;
assign te[1165] = 14;
assign s[1166] = 562751;
assign tm[1166] = 7681;
assign te[1166] = 14;
assign s[1167] = 566588;
assign tm[1167] = 7678;
assign te[1167] = 14;
assign s[1168] = 570424;
assign tm[1168] = 7675;
assign te[1168] = 14;
assign s[1169] = 574259;
assign tm[1169] = 7672;
assign te[1169] = 14;
assign s[1170] = 578092;
assign tm[1170] = 7668;
assign te[1170] = 14;
assign s[1171] = 581923;
assign tm[1171] = 7665;
assign te[1171] = 14;
assign s[1172] = 585753;
assign tm[1172] = 7662;
assign te[1172] = 14;
assign s[1173] = 589580;
assign tm[1173] = 7658;
assign te[1173] = 14;
assign s[1174] = 593407;
assign tm[1174] = 7655;
assign te[1174] = 14;
assign s[1175] = 597231;
assign tm[1175] = 7652;
assign te[1175] = 14;
assign s[1176] = 601054;
assign tm[1176] = 7649;
assign te[1176] = 14;
assign s[1177] = 604875;
assign tm[1177] = 7645;
assign te[1177] = 14;
assign s[1178] = 608695;
assign tm[1178] = 7642;
assign te[1178] = 14;
assign s[1179] = 612513;
assign tm[1179] = 7639;
assign te[1179] = 14;
assign s[1180] = 616330;
assign tm[1180] = 7636;
assign te[1180] = 14;
assign s[1181] = 620144;
assign tm[1181] = 7632;
assign te[1181] = 14;
assign s[1182] = 623958;
assign tm[1182] = 7629;
assign te[1182] = 14;
assign s[1183] = 627769;
assign tm[1183] = 7626;
assign te[1183] = 14;
assign s[1184] = 631579;
assign tm[1184] = 7623;
assign te[1184] = 14;
assign s[1185] = 635388;
assign tm[1185] = 7620;
assign te[1185] = 14;
assign s[1186] = 639195;
assign tm[1186] = 7616;
assign te[1186] = 14;
assign s[1187] = 643000;
assign tm[1187] = 7613;
assign te[1187] = 14;
assign s[1188] = 646803;
assign tm[1188] = 7610;
assign te[1188] = 14;
assign s[1189] = 650605;
assign tm[1189] = 7607;
assign te[1189] = 14;
assign s[1190] = 654406;
assign tm[1190] = 7603;
assign te[1190] = 14;
assign s[1191] = 658204;
assign tm[1191] = 7600;
assign te[1191] = 14;
assign s[1192] = 662002;
assign tm[1192] = 7597;
assign te[1192] = 14;
assign s[1193] = 665797;
assign tm[1193] = 7594;
assign te[1193] = 14;
assign s[1194] = 669591;
assign tm[1194] = 7591;
assign te[1194] = 14;
assign s[1195] = 673384;
assign tm[1195] = 7588;
assign te[1195] = 14;
assign s[1196] = 677175;
assign tm[1196] = 7584;
assign te[1196] = 14;
assign s[1197] = 680964;
assign tm[1197] = 7581;
assign te[1197] = 14;
assign s[1198] = 684751;
assign tm[1198] = 7578;
assign te[1198] = 14;
assign s[1199] = 688537;
assign tm[1199] = 7575;
assign te[1199] = 14;
assign s[1200] = 692322;
assign tm[1200] = 7572;
assign te[1200] = 14;
assign s[1201] = 696105;
assign tm[1201] = 7569;
assign te[1201] = 14;
assign s[1202] = 699887;
assign tm[1202] = 7565;
assign te[1202] = 14;
assign s[1203] = 703666;
assign tm[1203] = 7562;
assign te[1203] = 14;
assign s[1204] = 707444;
assign tm[1204] = 7559;
assign te[1204] = 14;
assign s[1205] = 711220;
assign tm[1205] = 7556;
assign te[1205] = 14;
assign s[1206] = 714996;
assign tm[1206] = 7553;
assign te[1206] = 14;
assign s[1207] = 718770;
assign tm[1207] = 7550;
assign te[1207] = 14;
assign s[1208] = 722542;
assign tm[1208] = 7547;
assign te[1208] = 14;
assign s[1209] = 726312;
assign tm[1209] = 7543;
assign te[1209] = 14;
assign s[1210] = 730080;
assign tm[1210] = 7540;
assign te[1210] = 14;
assign s[1211] = 733848;
assign tm[1211] = 7537;
assign te[1211] = 14;
assign s[1212] = 737614;
assign tm[1212] = 7534;
assign te[1212] = 14;
assign s[1213] = 741378;
assign tm[1213] = 7531;
assign te[1213] = 14;
assign s[1214] = 745141;
assign tm[1214] = 7528;
assign te[1214] = 14;
assign s[1215] = 748902;
assign tm[1215] = 7525;
assign te[1215] = 14;
assign s[1216] = 752661;
assign tm[1216] = 7522;
assign te[1216] = 14;
assign s[1217] = 756419;
assign tm[1217] = 7519;
assign te[1217] = 14;
assign s[1218] = 760175;
assign tm[1218] = 7515;
assign te[1218] = 14;
assign s[1219] = 763931;
assign tm[1219] = 7512;
assign te[1219] = 14;
assign s[1220] = 767684;
assign tm[1220] = 7509;
assign te[1220] = 14;
assign s[1221] = 771436;
assign tm[1221] = 7506;
assign te[1221] = 14;
assign s[1222] = 775186;
assign tm[1222] = 7503;
assign te[1222] = 14;
assign s[1223] = 778935;
assign tm[1223] = 7500;
assign te[1223] = 14;
assign s[1224] = 782682;
assign tm[1224] = 7497;
assign te[1224] = 14;
assign s[1225] = 786428;
assign tm[1225] = 7494;
assign te[1225] = 14;
assign s[1226] = 790172;
assign tm[1226] = 7491;
assign te[1226] = 14;
assign s[1227] = 793914;
assign tm[1227] = 7488;
assign te[1227] = 14;
assign s[1228] = 797655;
assign tm[1228] = 7485;
assign te[1228] = 14;
assign s[1229] = 801395;
assign tm[1229] = 7482;
assign te[1229] = 14;
assign s[1230] = 805133;
assign tm[1230] = 7479;
assign te[1230] = 14;
assign s[1231] = 808869;
assign tm[1231] = 7476;
assign te[1231] = 14;
assign s[1232] = 812604;
assign tm[1232] = 7473;
assign te[1232] = 14;
assign s[1233] = 816338;
assign tm[1233] = 7470;
assign te[1233] = 14;
assign s[1234] = 820070;
assign tm[1234] = 7466;
assign te[1234] = 14;
assign s[1235] = 823800;
assign tm[1235] = 7463;
assign te[1235] = 14;
assign s[1236] = 827529;
assign tm[1236] = 7460;
assign te[1236] = 14;
assign s[1237] = 831257;
assign tm[1237] = 7457;
assign te[1237] = 14;
assign s[1238] = 834983;
assign tm[1238] = 7454;
assign te[1238] = 14;
assign s[1239] = 838707;
assign tm[1239] = 7451;
assign te[1239] = 14;
assign s[1240] = 842430;
assign tm[1240] = 7448;
assign te[1240] = 14;
assign s[1241] = 846151;
assign tm[1241] = 7445;
assign te[1241] = 14;
assign s[1242] = 849872;
assign tm[1242] = 7442;
assign te[1242] = 14;
assign s[1243] = 853590;
assign tm[1243] = 7439;
assign te[1243] = 14;
assign s[1244] = 857307;
assign tm[1244] = 7436;
assign te[1244] = 14;
assign s[1245] = 861022;
assign tm[1245] = 7433;
assign te[1245] = 14;
assign s[1246] = 864736;
assign tm[1246] = 7430;
assign te[1246] = 14;
assign s[1247] = 868448;
assign tm[1247] = 7427;
assign te[1247] = 14;
assign s[1248] = 872160;
assign tm[1248] = 7424;
assign te[1248] = 14;
assign s[1249] = 875869;
assign tm[1249] = 7421;
assign te[1249] = 14;
assign s[1250] = 879578;
assign tm[1250] = 7418;
assign te[1250] = 14;
assign s[1251] = 883284;
assign tm[1251] = 7416;
assign te[1251] = 14;
assign s[1252] = 886989;
assign tm[1252] = 7413;
assign te[1252] = 14;
assign s[1253] = 890693;
assign tm[1253] = 7410;
assign te[1253] = 14;
assign s[1254] = 894395;
assign tm[1254] = 7407;
assign te[1254] = 14;
assign s[1255] = 898095;
assign tm[1255] = 7404;
assign te[1255] = 14;
assign s[1256] = 901794;
assign tm[1256] = 7401;
assign te[1256] = 14;
assign s[1257] = 905492;
assign tm[1257] = 7398;
assign te[1257] = 14;
assign s[1258] = 909188;
assign tm[1258] = 7395;
assign te[1258] = 14;
assign s[1259] = 912883;
assign tm[1259] = 7392;
assign te[1259] = 14;
assign s[1260] = 916577;
assign tm[1260] = 7389;
assign te[1260] = 14;
assign s[1261] = 920268;
assign tm[1261] = 7386;
assign te[1261] = 14;
assign s[1262] = 923958;
assign tm[1262] = 7383;
assign te[1262] = 14;
assign s[1263] = 927647;
assign tm[1263] = 7380;
assign te[1263] = 14;
assign s[1264] = 931334;
assign tm[1264] = 7377;
assign te[1264] = 14;
assign s[1265] = 935021;
assign tm[1265] = 7374;
assign te[1265] = 14;
assign s[1266] = 938705;
assign tm[1266] = 7371;
assign te[1266] = 14;
assign s[1267] = 942388;
assign tm[1267] = 7368;
assign te[1267] = 14;
assign s[1268] = 946070;
assign tm[1268] = 7366;
assign te[1268] = 14;
assign s[1269] = 949750;
assign tm[1269] = 7363;
assign te[1269] = 14;
assign s[1270] = 953428;
assign tm[1270] = 7360;
assign te[1270] = 14;
assign s[1271] = 957106;
assign tm[1271] = 7357;
assign te[1271] = 14;
assign s[1272] = 960782;
assign tm[1272] = 7354;
assign te[1272] = 14;
assign s[1273] = 964456;
assign tm[1273] = 7351;
assign te[1273] = 14;
assign s[1274] = 968129;
assign tm[1274] = 7348;
assign te[1274] = 14;
assign s[1275] = 971801;
assign tm[1275] = 7345;
assign te[1275] = 14;
assign s[1276] = 975470;
assign tm[1276] = 7342;
assign te[1276] = 14;
assign s[1277] = 979139;
assign tm[1277] = 7340;
assign te[1277] = 14;
assign s[1278] = 982807;
assign tm[1278] = 7337;
assign te[1278] = 14;
assign s[1279] = 986472;
assign tm[1279] = 7334;
assign te[1279] = 14;
assign s[1280] = 990136;
assign tm[1280] = 7331;
assign te[1280] = 14;
assign s[1281] = 993799;
assign tm[1281] = 7328;
assign te[1281] = 14;
assign s[1282] = 997461;
assign tm[1282] = 7325;
assign te[1282] = 14;
assign s[1283] = 1001121;
assign tm[1283] = 7322;
assign te[1283] = 14;
assign s[1284] = 1004779;
assign tm[1284] = 7319;
assign te[1284] = 14;
assign s[1285] = 1008437;
assign tm[1285] = 7317;
assign te[1285] = 14;
assign s[1286] = 1012092;
assign tm[1286] = 7314;
assign te[1286] = 14;
assign s[1287] = 1015746;
assign tm[1287] = 7311;
assign te[1287] = 14;
assign s[1288] = 1019400;
assign tm[1288] = 7308;
assign te[1288] = 14;
assign s[1289] = 1023051;
assign tm[1289] = 7305;
assign te[1289] = 14;
assign s[1290] = 1026701;
assign tm[1290] = 7302;
assign te[1290] = 14;
assign s[1291] = 1030350;
assign tm[1291] = 7300;
assign te[1291] = 14;
assign s[1292] = 1033997;
assign tm[1292] = 7297;
assign te[1292] = 14;
assign s[1293] = 1037643;
assign tm[1293] = 7294;
assign te[1293] = 14;
assign s[1294] = 1041287;
assign tm[1294] = 7291;
assign te[1294] = 14;
assign s[1295] = 1044930;
assign tm[1295] = 7288;
assign te[1295] = 14;
assign s[1296] = 1048571;
assign tm[1296] = 7285;
assign te[1296] = 14;
assign s[1297] = 1052211;
assign tm[1297] = 7283;
assign te[1297] = 14;
assign s[1298] = 1055851;
assign tm[1298] = 7280;
assign te[1298] = 14;
assign s[1299] = 1059488;
assign tm[1299] = 7277;
assign te[1299] = 14;
assign s[1300] = 1063123;
assign tm[1300] = 7274;
assign te[1300] = 14;
assign s[1301] = 1066759;
assign tm[1301] = 7271;
assign te[1301] = 14;
assign s[1302] = 1070392;
assign tm[1302] = 7269;
assign te[1302] = 14;
assign s[1303] = 1074023;
assign tm[1303] = 7266;
assign te[1303] = 14;
assign s[1304] = 1077654;
assign tm[1304] = 7263;
assign te[1304] = 14;
assign s[1305] = 1081283;
assign tm[1305] = 7260;
assign te[1305] = 14;
assign s[1306] = 1084911;
assign tm[1306] = 7258;
assign te[1306] = 14;
assign s[1307] = 1088537;
assign tm[1307] = 7255;
assign te[1307] = 14;
assign s[1308] = 1092161;
assign tm[1308] = 7252;
assign te[1308] = 14;
assign s[1309] = 1095785;
assign tm[1309] = 7249;
assign te[1309] = 14;
assign s[1310] = 1099407;
assign tm[1310] = 7246;
assign te[1310] = 14;
assign s[1311] = 1103028;
assign tm[1311] = 7244;
assign te[1311] = 14;
assign s[1312] = 1106647;
assign tm[1312] = 7241;
assign te[1312] = 14;
assign s[1313] = 1110265;
assign tm[1313] = 7238;
assign te[1313] = 14;
assign s[1314] = 1113882;
assign tm[1314] = 7235;
assign te[1314] = 14;
assign s[1315] = 1117497;
assign tm[1315] = 7233;
assign te[1315] = 14;
assign s[1316] = 1121110;
assign tm[1316] = 7230;
assign te[1316] = 14;
assign s[1317] = 1124723;
assign tm[1317] = 7227;
assign te[1317] = 14;
assign s[1318] = 1128334;
assign tm[1318] = 7224;
assign te[1318] = 14;
assign s[1319] = 1131944;
assign tm[1319] = 7222;
assign te[1319] = 14;
assign s[1320] = 1135552;
assign tm[1320] = 7219;
assign te[1320] = 14;
assign s[1321] = 1139159;
assign tm[1321] = 7216;
assign te[1321] = 14;
assign s[1322] = 1142765;
assign tm[1322] = 7213;
assign te[1322] = 14;
assign s[1323] = 1146369;
assign tm[1323] = 7211;
assign te[1323] = 14;
assign s[1324] = 1149971;
assign tm[1324] = 7208;
assign te[1324] = 14;
assign s[1325] = 1153573;
assign tm[1325] = 7205;
assign te[1325] = 14;
assign s[1326] = 1157173;
assign tm[1326] = 7203;
assign te[1326] = 14;
assign s[1327] = 1160772;
assign tm[1327] = 7200;
assign te[1327] = 14;
assign s[1328] = 1164369;
assign tm[1328] = 7197;
assign te[1328] = 14;
assign s[1329] = 1167965;
assign tm[1329] = 7194;
assign te[1329] = 14;
assign s[1330] = 1171560;
assign tm[1330] = 7192;
assign te[1330] = 14;
assign s[1331] = 1175153;
assign tm[1331] = 7189;
assign te[1331] = 14;
assign s[1332] = 1178746;
assign tm[1332] = 7186;
assign te[1332] = 14;
assign s[1333] = 1182336;
assign tm[1333] = 7184;
assign te[1333] = 14;
assign s[1334] = 1185926;
assign tm[1334] = 7181;
assign te[1334] = 14;
assign s[1335] = 1189513;
assign tm[1335] = 7178;
assign te[1335] = 14;
assign s[1336] = 1193100;
assign tm[1336] = 7175;
assign te[1336] = 14;
assign s[1337] = 1196685;
assign tm[1337] = 7173;
assign te[1337] = 14;
assign s[1338] = 1200270;
assign tm[1338] = 7170;
assign te[1338] = 14;
assign s[1339] = 1203852;
assign tm[1339] = 7167;
assign te[1339] = 14;
assign s[1340] = 1207434;
assign tm[1340] = 7165;
assign te[1340] = 14;
assign s[1341] = 1211013;
assign tm[1341] = 7162;
assign te[1341] = 14;
assign s[1342] = 1214592;
assign tm[1342] = 7159;
assign te[1342] = 14;
assign s[1343] = 1218170;
assign tm[1343] = 7157;
assign te[1343] = 14;
assign s[1344] = 1221746;
assign tm[1344] = 7154;
assign te[1344] = 14;
assign s[1345] = 1225320;
assign tm[1345] = 7151;
assign te[1345] = 14;
assign s[1346] = 1228893;
assign tm[1346] = 7149;
assign te[1346] = 14;
assign s[1347] = 1232465;
assign tm[1347] = 7146;
assign te[1347] = 14;
assign s[1348] = 1236036;
assign tm[1348] = 7143;
assign te[1348] = 14;
assign s[1349] = 1239605;
assign tm[1349] = 7141;
assign te[1349] = 14;
assign s[1350] = 1243173;
assign tm[1350] = 7138;
assign te[1350] = 14;
assign s[1351] = 1246740;
assign tm[1351] = 7135;
assign te[1351] = 14;
assign s[1352] = 1250305;
assign tm[1352] = 7133;
assign te[1352] = 14;
assign s[1353] = 1253870;
assign tm[1353] = 7130;
assign te[1353] = 14;
assign s[1354] = 1257432;
assign tm[1354] = 7128;
assign te[1354] = 14;
assign s[1355] = 1260993;
assign tm[1355] = 7125;
assign te[1355] = 14;
assign s[1356] = 1264553;
assign tm[1356] = 7122;
assign te[1356] = 14;
assign s[1357] = 1268113;
assign tm[1357] = 7120;
assign te[1357] = 14;
assign s[1358] = 1271670;
assign tm[1358] = 7117;
assign te[1358] = 14;
assign s[1359] = 1275226;
assign tm[1359] = 7114;
assign te[1359] = 14;
assign s[1360] = 1278780;
assign tm[1360] = 7112;
assign te[1360] = 14;
assign s[1361] = 1282334;
assign tm[1361] = 7109;
assign te[1361] = 14;
assign s[1362] = 1285886;
assign tm[1362] = 7107;
assign te[1362] = 14;
assign s[1363] = 1289437;
assign tm[1363] = 7104;
assign te[1363] = 14;
assign s[1364] = 1292987;
assign tm[1364] = 7101;
assign te[1364] = 14;
assign s[1365] = 1296535;
assign tm[1365] = 7099;
assign te[1365] = 14;
assign s[1366] = 1300082;
assign tm[1366] = 7096;
assign te[1366] = 14;
assign s[1367] = 1303628;
assign tm[1367] = 7094;
assign te[1367] = 14;
assign s[1368] = 1307173;
assign tm[1368] = 7091;
assign te[1368] = 14;
assign s[1369] = 1310716;
assign tm[1369] = 7088;
assign te[1369] = 14;
assign s[1370] = 1314258;
assign tm[1370] = 7086;
assign te[1370] = 14;
assign s[1371] = 1317798;
assign tm[1371] = 7083;
assign te[1371] = 14;
assign s[1372] = 1321337;
assign tm[1372] = 7081;
assign te[1372] = 14;
assign s[1373] = 1324875;
assign tm[1373] = 7078;
assign te[1373] = 14;
assign s[1374] = 1328412;
assign tm[1374] = 7075;
assign te[1374] = 14;
assign s[1375] = 1331948;
assign tm[1375] = 7073;
assign te[1375] = 14;
assign s[1376] = 1335481;
assign tm[1376] = 7070;
assign te[1376] = 14;
assign s[1377] = 1339014;
assign tm[1377] = 7068;
assign te[1377] = 14;
assign s[1378] = 1342546;
assign tm[1378] = 7065;
assign te[1378] = 14;
assign s[1379] = 1346076;
assign tm[1379] = 7063;
assign te[1379] = 14;
assign s[1380] = 1349605;
assign tm[1380] = 7060;
assign te[1380] = 14;
assign s[1381] = 1353133;
assign tm[1381] = 7057;
assign te[1381] = 14;
assign s[1382] = 1356659;
assign tm[1382] = 7055;
assign te[1382] = 14;
assign s[1383] = 1360184;
assign tm[1383] = 7052;
assign te[1383] = 14;
assign s[1384] = 1363708;
assign tm[1384] = 7050;
assign te[1384] = 14;
assign s[1385] = 1367230;
assign tm[1385] = 7047;
assign te[1385] = 14;
assign s[1386] = 1370752;
assign tm[1386] = 7045;
assign te[1386] = 14;
assign s[1387] = 1374272;
assign tm[1387] = 7042;
assign te[1387] = 14;
assign s[1388] = 1377791;
assign tm[1388] = 7040;
assign te[1388] = 14;
assign s[1389] = 1381308;
assign tm[1389] = 7037;
assign te[1389] = 14;
assign s[1390] = 1384824;
assign tm[1390] = 7035;
assign te[1390] = 14;
assign s[1391] = 1388340;
assign tm[1391] = 7032;
assign te[1391] = 14;
assign s[1392] = 1391853;
assign tm[1392] = 7029;
assign te[1392] = 14;
assign s[1393] = 1395366;
assign tm[1393] = 7027;
assign te[1393] = 14;
assign s[1394] = 1398877;
assign tm[1394] = 7024;
assign te[1394] = 14;
assign s[1395] = 1402387;
assign tm[1395] = 7022;
assign te[1395] = 14;
assign s[1396] = 1405896;
assign tm[1396] = 7019;
assign te[1396] = 14;
assign s[1397] = 1409403;
assign tm[1397] = 7017;
assign te[1397] = 14;
assign s[1398] = 1412909;
assign tm[1398] = 7014;
assign te[1398] = 14;
assign s[1399] = 1416414;
assign tm[1399] = 7012;
assign te[1399] = 14;
assign s[1400] = 1419918;
assign tm[1400] = 7009;
assign te[1400] = 14;
assign s[1401] = 1423420;
assign tm[1401] = 7007;
assign te[1401] = 14;
assign s[1402] = 1426921;
assign tm[1402] = 7004;
assign te[1402] = 14;
assign s[1403] = 1430421;
assign tm[1403] = 7002;
assign te[1403] = 14;
assign s[1404] = 1433920;
assign tm[1404] = 6999;
assign te[1404] = 14;
assign s[1405] = 1437418;
assign tm[1405] = 6997;
assign te[1405] = 14;
assign s[1406] = 1440914;
assign tm[1406] = 6994;
assign te[1406] = 14;
assign s[1407] = 1444409;
assign tm[1407] = 6992;
assign te[1407] = 14;
assign s[1408] = 1447902;
assign tm[1408] = 6989;
assign te[1408] = 14;
assign s[1409] = 1451395;
assign tm[1409] = 6987;
assign te[1409] = 14;
assign s[1410] = 1454886;
assign tm[1410] = 6984;
assign te[1410] = 14;
assign s[1411] = 1458376;
assign tm[1411] = 6982;
assign te[1411] = 14;
assign s[1412] = 1461865;
assign tm[1412] = 6979;
assign te[1412] = 14;
assign s[1413] = 1465352;
assign tm[1413] = 6977;
assign te[1413] = 14;
assign s[1414] = 1468838;
assign tm[1414] = 6975;
assign te[1414] = 14;
assign s[1415] = 1472324;
assign tm[1415] = 6972;
assign te[1415] = 14;
assign s[1416] = 1475807;
assign tm[1416] = 6970;
assign te[1416] = 14;
assign s[1417] = 1479290;
assign tm[1417] = 6967;
assign te[1417] = 14;
assign s[1418] = 1482771;
assign tm[1418] = 6965;
assign te[1418] = 14;
assign s[1419] = 1486251;
assign tm[1419] = 6962;
assign te[1419] = 14;
assign s[1420] = 1489730;
assign tm[1420] = 6960;
assign te[1420] = 14;
assign s[1421] = 1493208;
assign tm[1421] = 6957;
assign te[1421] = 14;
assign s[1422] = 1496684;
assign tm[1422] = 6955;
assign te[1422] = 14;
assign s[1423] = 1500160;
assign tm[1423] = 6952;
assign te[1423] = 14;
assign s[1424] = 1503634;
assign tm[1424] = 6950;
assign te[1424] = 14;
assign s[1425] = 1507107;
assign tm[1425] = 6948;
assign te[1425] = 14;
assign s[1426] = 1510578;
assign tm[1426] = 6945;
assign te[1426] = 14;
assign s[1427] = 1514048;
assign tm[1427] = 6943;
assign te[1427] = 14;
assign s[1428] = 1517518;
assign tm[1428] = 6940;
assign te[1428] = 14;
assign s[1429] = 1520986;
assign tm[1429] = 6938;
assign te[1429] = 14;
assign s[1430] = 1524453;
assign tm[1430] = 6935;
assign te[1430] = 14;
assign s[1431] = 1527918;
assign tm[1431] = 6933;
assign te[1431] = 14;
assign s[1432] = 1531382;
assign tm[1432] = 6930;
assign te[1432] = 14;
assign s[1433] = 1534845;
assign tm[1433] = 6928;
assign te[1433] = 14;
assign s[1434] = 1538307;
assign tm[1434] = 6926;
assign te[1434] = 14;
assign s[1435] = 1541768;
assign tm[1435] = 6923;
assign te[1435] = 14;
assign s[1436] = 1545227;
assign tm[1436] = 6921;
assign te[1436] = 14;
assign s[1437] = 1548685;
assign tm[1437] = 6918;
assign te[1437] = 14;
assign s[1438] = 1552142;
assign tm[1438] = 6916;
assign te[1438] = 14;
assign s[1439] = 1555599;
assign tm[1439] = 6914;
assign te[1439] = 14;
assign s[1440] = 1559053;
assign tm[1440] = 6911;
assign te[1440] = 14;
assign s[1441] = 1562506;
assign tm[1441] = 6909;
assign te[1441] = 14;
assign s[1442] = 1565958;
assign tm[1442] = 6906;
assign te[1442] = 14;
assign s[1443] = 1569410;
assign tm[1443] = 6904;
assign te[1443] = 14;
assign s[1444] = 1572859;
assign tm[1444] = 6902;
assign te[1444] = 14;
assign s[1445] = 1576308;
assign tm[1445] = 6899;
assign te[1445] = 14;
assign s[1446] = 1579756;
assign tm[1446] = 6897;
assign te[1446] = 14;
assign s[1447] = 1583202;
assign tm[1447] = 6894;
assign te[1447] = 14;
assign s[1448] = 1586647;
assign tm[1448] = 6892;
assign te[1448] = 14;
assign s[1449] = 1590090;
assign tm[1449] = 6890;
assign te[1449] = 14;
assign s[1450] = 1593534;
assign tm[1450] = 6887;
assign te[1450] = 14;
assign s[1451] = 1596975;
assign tm[1451] = 6885;
assign te[1451] = 14;
assign s[1452] = 1600416;
assign tm[1452] = 6883;
assign te[1452] = 14;
assign s[1453] = 1603854;
assign tm[1453] = 6880;
assign te[1453] = 14;
assign s[1454] = 1607293;
assign tm[1454] = 6878;
assign te[1454] = 14;
assign s[1455] = 1610729;
assign tm[1455] = 6875;
assign te[1455] = 14;
assign s[1456] = 1614165;
assign tm[1456] = 6873;
assign te[1456] = 14;
assign s[1457] = 1617599;
assign tm[1457] = 6871;
assign te[1457] = 14;
assign s[1458] = 1621033;
assign tm[1458] = 6868;
assign te[1458] = 14;
assign s[1459] = 1624465;
assign tm[1459] = 6866;
assign te[1459] = 14;
assign s[1460] = 1627896;
assign tm[1460] = 6864;
assign te[1460] = 14;
assign s[1461] = 1631325;
assign tm[1461] = 6861;
assign te[1461] = 14;
assign s[1462] = 1634754;
assign tm[1462] = 6859;
assign te[1462] = 14;
assign s[1463] = 1638182;
assign tm[1463] = 6857;
assign te[1463] = 14;
assign s[1464] = 1641607;
assign tm[1464] = 6854;
assign te[1464] = 14;
assign s[1465] = 1645033;
assign tm[1465] = 6852;
assign te[1465] = 14;
assign s[1466] = 1648457;
assign tm[1466] = 6850;
assign te[1466] = 14;
assign s[1467] = 1651879;
assign tm[1467] = 6847;
assign te[1467] = 14;
assign s[1468] = 1655301;
assign tm[1468] = 6845;
assign te[1468] = 14;
assign s[1469] = 1658721;
assign tm[1469] = 6843;
assign te[1469] = 14;
assign s[1470] = 1662140;
assign tm[1470] = 6840;
assign te[1470] = 14;
assign s[1471] = 1665558;
assign tm[1471] = 6838;
assign te[1471] = 14;
assign s[1472] = 1668975;
assign tm[1472] = 6836;
assign te[1472] = 14;
assign s[1473] = 1672391;
assign tm[1473] = 6833;
assign te[1473] = 14;
assign s[1474] = 1675806;
assign tm[1474] = 6831;
assign te[1474] = 14;
assign s[1475] = 1679219;
assign tm[1475] = 6829;
assign te[1475] = 14;
assign s[1476] = 1682631;
assign tm[1476] = 6826;
assign te[1476] = 14;
assign s[1477] = 1686042;
assign tm[1477] = 6824;
assign te[1477] = 14;
assign s[1478] = 1689452;
assign tm[1478] = 6822;
assign te[1478] = 14;
assign s[1479] = 1692861;
assign tm[1479] = 6819;
assign te[1479] = 14;
assign s[1480] = 1696269;
assign tm[1480] = 6817;
assign te[1480] = 14;
assign s[1481] = 1699675;
assign tm[1481] = 6815;
assign te[1481] = 14;
assign s[1482] = 1703081;
assign tm[1482] = 6812;
assign te[1482] = 14;
assign s[1483] = 1706485;
assign tm[1483] = 6810;
assign te[1483] = 14;
assign s[1484] = 1709888;
assign tm[1484] = 6808;
assign te[1484] = 14;
assign s[1485] = 1713290;
assign tm[1485] = 6806;
assign te[1485] = 14;
assign s[1486] = 1716690;
assign tm[1486] = 6803;
assign te[1486] = 14;
assign s[1487] = 1720090;
assign tm[1487] = 6801;
assign te[1487] = 14;
assign s[1488] = 1723488;
assign tm[1488] = 6799;
assign te[1488] = 14;
assign s[1489] = 1726886;
assign tm[1489] = 6796;
assign te[1489] = 14;
assign s[1490] = 1730282;
assign tm[1490] = 6794;
assign te[1490] = 14;
assign s[1491] = 1733677;
assign tm[1491] = 6792;
assign te[1491] = 14;
assign s[1492] = 1737070;
assign tm[1492] = 6790;
assign te[1492] = 14;
assign s[1493] = 1740463;
assign tm[1493] = 6787;
assign te[1493] = 14;
assign s[1494] = 1743855;
assign tm[1494] = 6785;
assign te[1494] = 14;
assign s[1495] = 1747246;
assign tm[1495] = 6783;
assign te[1495] = 14;
assign s[1496] = 1750635;
assign tm[1496] = 6780;
assign te[1496] = 14;
assign s[1497] = 1754023;
assign tm[1497] = 6778;
assign te[1497] = 14;
assign s[1498] = 1757410;
assign tm[1498] = 6776;
assign te[1498] = 14;
assign s[1499] = 1760796;
assign tm[1499] = 6774;
assign te[1499] = 14;
assign s[1500] = 1764181;
assign tm[1500] = 6771;
assign te[1500] = 14;
assign s[1501] = 1767565;
assign tm[1501] = 6769;
assign te[1501] = 14;
assign s[1502] = 1770947;
assign tm[1502] = 6767;
assign te[1502] = 14;
assign s[1503] = 1774328;
assign tm[1503] = 6765;
assign te[1503] = 14;
assign s[1504] = 1777709;
assign tm[1504] = 6762;
assign te[1504] = 14;
assign s[1505] = 1781088;
assign tm[1505] = 6760;
assign te[1505] = 14;
assign s[1506] = 1784467;
assign tm[1506] = 6758;
assign te[1506] = 14;
assign s[1507] = 1787844;
assign tm[1507] = 6756;
assign te[1507] = 14;
assign s[1508] = 1791219;
assign tm[1508] = 6753;
assign te[1508] = 14;
assign s[1509] = 1794594;
assign tm[1509] = 6751;
assign te[1509] = 14;
assign s[1510] = 1797967;
assign tm[1510] = 6749;
assign te[1510] = 14;
assign s[1511] = 1801340;
assign tm[1511] = 6747;
assign te[1511] = 14;
assign s[1512] = 1804711;
assign tm[1512] = 6744;
assign te[1512] = 14;
assign s[1513] = 1808081;
assign tm[1513] = 6742;
assign te[1513] = 14;
assign s[1514] = 1811450;
assign tm[1514] = 6740;
assign te[1514] = 14;
assign s[1515] = 1814819;
assign tm[1515] = 6738;
assign te[1515] = 14;
assign s[1516] = 1818186;
assign tm[1516] = 6736;
assign te[1516] = 14;
assign s[1517] = 1821552;
assign tm[1517] = 6733;
assign te[1517] = 14;
assign s[1518] = 1824916;
assign tm[1518] = 6731;
assign te[1518] = 14;
assign s[1519] = 1828280;
assign tm[1519] = 6729;
assign te[1519] = 14;
assign s[1520] = 1831643;
assign tm[1520] = 6727;
assign te[1520] = 14;
assign s[1521] = 1835003;
assign tm[1521] = 6724;
assign te[1521] = 14;
assign s[1522] = 1838364;
assign tm[1522] = 6722;
assign te[1522] = 14;
assign s[1523] = 1841723;
assign tm[1523] = 6720;
assign te[1523] = 14;
assign s[1524] = 1845082;
assign tm[1524] = 6718;
assign te[1524] = 14;
assign s[1525] = 1848438;
assign tm[1525] = 6716;
assign te[1525] = 14;
assign s[1526] = 1851794;
assign tm[1526] = 6713;
assign te[1526] = 14;
assign s[1527] = 1855148;
assign tm[1527] = 6711;
assign te[1527] = 14;
assign s[1528] = 1858502;
assign tm[1528] = 6709;
assign te[1528] = 14;
assign s[1529] = 1861855;
assign tm[1529] = 6707;
assign te[1529] = 14;
assign s[1530] = 1865206;
assign tm[1530] = 6705;
assign te[1530] = 14;
assign s[1531] = 1868557;
assign tm[1531] = 6702;
assign te[1531] = 14;
assign s[1532] = 1871906;
assign tm[1532] = 6700;
assign te[1532] = 14;
assign s[1533] = 1875254;
assign tm[1533] = 6698;
assign te[1533] = 14;
assign s[1534] = 1878601;
assign tm[1534] = 6696;
assign te[1534] = 14;
assign s[1535] = 1881948;
assign tm[1535] = 6694;
assign te[1535] = 14;
assign s[1536] = 1885292;
assign tm[1536] = 6692;
assign te[1536] = 14;
assign s[1537] = 1888636;
assign tm[1537] = 6689;
assign te[1537] = 14;
assign s[1538] = 1891979;
assign tm[1538] = 6687;
assign te[1538] = 14;
assign s[1539] = 1895320;
assign tm[1539] = 6685;
assign te[1539] = 14;
assign s[1540] = 1898661;
assign tm[1540] = 6683;
assign te[1540] = 14;
assign s[1541] = 1902000;
assign tm[1541] = 6681;
assign te[1541] = 14;
assign s[1542] = 1905339;
assign tm[1542] = 6678;
assign te[1542] = 14;
assign s[1543] = 1908676;
assign tm[1543] = 6676;
assign te[1543] = 14;
assign s[1544] = 1912012;
assign tm[1544] = 6674;
assign te[1544] = 14;
assign s[1545] = 1915348;
assign tm[1545] = 6672;
assign te[1545] = 14;
assign s[1546] = 1918682;
assign tm[1546] = 6670;
assign te[1546] = 14;
assign s[1547] = 1922014;
assign tm[1547] = 6668;
assign te[1547] = 14;
assign s[1548] = 1925347;
assign tm[1548] = 6665;
assign te[1548] = 14;
assign s[1549] = 1928677;
assign tm[1549] = 6663;
assign te[1549] = 14;
assign s[1550] = 1932007;
assign tm[1550] = 6661;
assign te[1550] = 14;
assign s[1551] = 1935336;
assign tm[1551] = 6659;
assign te[1551] = 14;
assign s[1552] = 1938663;
assign tm[1552] = 6657;
assign te[1552] = 14;
assign s[1553] = 1941990;
assign tm[1553] = 6655;
assign te[1553] = 14;
assign s[1554] = 1945316;
assign tm[1554] = 6653;
assign te[1554] = 14;
assign s[1555] = 1948640;
assign tm[1555] = 6650;
assign te[1555] = 14;
assign s[1556] = 1951963;
assign tm[1556] = 6648;
assign te[1556] = 14;
assign s[1557] = 1955286;
assign tm[1557] = 6646;
assign te[1557] = 14;
assign s[1558] = 1958607;
assign tm[1558] = 6644;
assign te[1558] = 14;
assign s[1559] = 1961927;
assign tm[1559] = 6642;
assign te[1559] = 14;
assign s[1560] = 1965246;
assign tm[1560] = 6640;
assign te[1560] = 14;
assign s[1561] = 1968564;
assign tm[1561] = 6638;
assign te[1561] = 14;
assign s[1562] = 1971881;
assign tm[1562] = 6636;
assign te[1562] = 14;
assign s[1563] = 1975197;
assign tm[1563] = 6633;
assign te[1563] = 14;
assign s[1564] = 1978512;
assign tm[1564] = 6631;
assign te[1564] = 14;
assign s[1565] = 1981826;
assign tm[1565] = 6629;
assign te[1565] = 14;
assign s[1566] = 1985138;
assign tm[1566] = 6627;
assign te[1566] = 14;
assign s[1567] = 1988450;
assign tm[1567] = 6625;
assign te[1567] = 14;
assign s[1568] = 1991760;
assign tm[1568] = 6623;
assign te[1568] = 14;
assign s[1569] = 1995070;
assign tm[1569] = 6621;
assign te[1569] = 14;
assign s[1570] = 1998379;
assign tm[1570] = 6619;
assign te[1570] = 14;
assign s[1571] = 2001686;
assign tm[1571] = 6616;
assign te[1571] = 14;
assign s[1572] = 2004992;
assign tm[1572] = 6614;
assign te[1572] = 14;
assign s[1573] = 2008298;
assign tm[1573] = 6612;
assign te[1573] = 14;
assign s[1574] = 2011602;
assign tm[1574] = 6610;
assign te[1574] = 14;
assign s[1575] = 2014905;
assign tm[1575] = 6608;
assign te[1575] = 14;
assign s[1576] = 2018207;
assign tm[1576] = 6606;
assign te[1576] = 14;
assign s[1577] = 2021509;
assign tm[1577] = 6604;
assign te[1577] = 14;
assign s[1578] = 2024808;
assign tm[1578] = 6602;
assign te[1578] = 14;
assign s[1579] = 2028108;
assign tm[1579] = 6600;
assign te[1579] = 14;
assign s[1580] = 2031405;
assign tm[1580] = 6598;
assign te[1580] = 14;
assign s[1581] = 2034703;
assign tm[1581] = 6595;
assign te[1581] = 14;
assign s[1582] = 2037998;
assign tm[1582] = 6593;
assign te[1582] = 14;
assign s[1583] = 2041294;
assign tm[1583] = 6591;
assign te[1583] = 14;
assign s[1584] = 2044587;
assign tm[1584] = 6589;
assign te[1584] = 14;
assign s[1585] = 2047880;
assign tm[1585] = 6587;
assign te[1585] = 14;
assign s[1586] = 2051171;
assign tm[1586] = 6585;
assign te[1586] = 14;
assign s[1587] = 2054463;
assign tm[1587] = 6583;
assign te[1587] = 14;
assign s[1588] = 2057752;
assign tm[1588] = 6581;
assign te[1588] = 14;
assign s[1589] = 2061041;
assign tm[1589] = 6579;
assign te[1589] = 14;
assign s[1590] = 2064329;
assign tm[1590] = 6577;
assign te[1590] = 14;
assign s[1591] = 2067615;
assign tm[1591] = 6575;
assign te[1591] = 14;
assign s[1592] = 2070901;
assign tm[1592] = 6573;
assign te[1592] = 14;
assign s[1593] = 2074184;
assign tm[1593] = 6571;
assign te[1593] = 14;
assign s[1594] = 2077469;
assign tm[1594] = 6569;
assign te[1594] = 14;
assign s[1595] = 2080751;
assign tm[1595] = 6566;
assign te[1595] = 14;
assign s[1596] = 2084032;
assign tm[1596] = 6564;
assign te[1596] = 14;
assign s[1597] = 2087313;
assign tm[1597] = 6562;
assign te[1597] = 14;
assign s[1598] = 2090592;
assign tm[1598] = 6560;
assign te[1598] = 14;
assign s[1599] = 2093870;
assign tm[1599] = 6558;
assign te[1599] = 14;
assign s[1600] = 2097147;
assign tm[1600] = 6556;
assign te[1600] = 14;
assign s[1601] = 2100423;
assign tm[1601] = 6554;
assign te[1601] = 14;
assign s[1602] = 2103699;
assign tm[1602] = 6552;
assign te[1602] = 14;
assign s[1603] = 2106973;
assign tm[1603] = 6550;
assign te[1603] = 14;
assign s[1604] = 2110246;
assign tm[1604] = 6548;
assign te[1604] = 14;
assign s[1605] = 2113519;
assign tm[1605] = 6546;
assign te[1605] = 14;
assign s[1606] = 2116790;
assign tm[1606] = 6544;
assign te[1606] = 14;
assign s[1607] = 2120061;
assign tm[1607] = 6542;
assign te[1607] = 14;
assign s[1608] = 2123329;
assign tm[1608] = 6540;
assign te[1608] = 14;
assign s[1609] = 2126598;
assign tm[1609] = 6538;
assign te[1609] = 14;
assign s[1610] = 2129865;
assign tm[1610] = 6536;
assign te[1610] = 14;
assign s[1611] = 2133131;
assign tm[1611] = 6534;
assign te[1611] = 14;
assign s[1612] = 2136396;
assign tm[1612] = 6532;
assign te[1612] = 14;
assign s[1613] = 2139659;
assign tm[1613] = 6530;
assign te[1613] = 14;
assign s[1614] = 2142923;
assign tm[1614] = 6528;
assign te[1614] = 14;
assign s[1615] = 2146185;
assign tm[1615] = 6526;
assign te[1615] = 14;
assign s[1616] = 2149446;
assign tm[1616] = 6524;
assign te[1616] = 14;
assign s[1617] = 2152706;
assign tm[1617] = 6522;
assign te[1617] = 14;
assign s[1618] = 2155965;
assign tm[1618] = 6520;
assign te[1618] = 14;
assign s[1619] = 2159223;
assign tm[1619] = 6518;
assign te[1619] = 14;
assign s[1620] = 2162480;
assign tm[1620] = 6516;
assign te[1620] = 14;
assign s[1621] = 2165736;
assign tm[1621] = 6514;
assign te[1621] = 14;
assign s[1622] = 2168991;
assign tm[1622] = 6512;
assign te[1622] = 14;
assign s[1623] = 2172245;
assign tm[1623] = 6510;
assign te[1623] = 14;
assign s[1624] = 2175498;
assign tm[1624] = 6507;
assign te[1624] = 14;
assign s[1625] = 2178750;
assign tm[1625] = 6505;
assign te[1625] = 14;
assign s[1626] = 2182001;
assign tm[1626] = 6503;
assign te[1626] = 14;
assign s[1627] = 2185251;
assign tm[1627] = 6501;
assign te[1627] = 14;
assign s[1628] = 2188500;
assign tm[1628] = 6499;
assign te[1628] = 14;
assign s[1629] = 2191748;
assign tm[1629] = 6497;
assign te[1629] = 14;
assign s[1630] = 2194995;
assign tm[1630] = 6495;
assign te[1630] = 14;
assign s[1631] = 2198241;
assign tm[1631] = 6494;
assign te[1631] = 14;
assign s[1632] = 2201486;
assign tm[1632] = 6492;
assign te[1632] = 14;
assign s[1633] = 2204730;
assign tm[1633] = 6490;
assign te[1633] = 14;
assign s[1634] = 2207973;
assign tm[1634] = 6488;
assign te[1634] = 14;
assign s[1635] = 2211215;
assign tm[1635] = 6486;
assign te[1635] = 14;
assign s[1636] = 2214456;
assign tm[1636] = 6484;
assign te[1636] = 14;
assign s[1637] = 2217696;
assign tm[1637] = 6482;
assign te[1637] = 14;
assign s[1638] = 2220936;
assign tm[1638] = 6480;
assign te[1638] = 14;
assign s[1639] = 2224174;
assign tm[1639] = 6478;
assign te[1639] = 14;
assign s[1640] = 2227410;
assign tm[1640] = 6476;
assign te[1640] = 14;
assign s[1641] = 2230646;
assign tm[1641] = 6474;
assign te[1641] = 14;
assign s[1642] = 2233882;
assign tm[1642] = 6472;
assign te[1642] = 14;
assign s[1643] = 2237116;
assign tm[1643] = 6470;
assign te[1643] = 14;
assign s[1644] = 2240349;
assign tm[1644] = 6468;
assign te[1644] = 14;
assign s[1645] = 2243581;
assign tm[1645] = 6466;
assign te[1645] = 14;
assign s[1646] = 2246813;
assign tm[1646] = 6464;
assign te[1646] = 14;
assign s[1647] = 2250043;
assign tm[1647] = 6462;
assign te[1647] = 14;
assign s[1648] = 2253272;
assign tm[1648] = 6460;
assign te[1648] = 14;
assign s[1649] = 2256500;
assign tm[1649] = 6458;
assign te[1649] = 14;
assign s[1650] = 2259727;
assign tm[1650] = 6456;
assign te[1650] = 14;
assign s[1651] = 2262953;
assign tm[1651] = 6454;
assign te[1651] = 14;
assign s[1652] = 2266179;
assign tm[1652] = 6452;
assign te[1652] = 14;
assign s[1653] = 2269403;
assign tm[1653] = 6450;
assign te[1653] = 14;
assign s[1654] = 2272626;
assign tm[1654] = 6448;
assign te[1654] = 14;
assign s[1655] = 2275849;
assign tm[1655] = 6446;
assign te[1655] = 14;
assign s[1656] = 2279070;
assign tm[1656] = 6444;
assign te[1656] = 14;
assign s[1657] = 2282291;
assign tm[1657] = 6442;
assign te[1657] = 14;
assign s[1658] = 2285510;
assign tm[1658] = 6440;
assign te[1658] = 14;
assign s[1659] = 2288729;
assign tm[1659] = 6438;
assign te[1659] = 14;
assign s[1660] = 2291946;
assign tm[1660] = 6436;
assign te[1660] = 14;
assign s[1661] = 2295163;
assign tm[1661] = 6435;
assign te[1661] = 14;
assign s[1662] = 2298378;
assign tm[1662] = 6433;
assign te[1662] = 14;
assign s[1663] = 2301593;
assign tm[1663] = 6431;
assign te[1663] = 14;
assign s[1664] = 2304807;
assign tm[1664] = 6429;
assign te[1664] = 14;
assign s[1665] = 2308019;
assign tm[1665] = 6427;
assign te[1665] = 14;
assign s[1666] = 2311231;
assign tm[1666] = 6425;
assign te[1666] = 14;
assign s[1667] = 2314442;
assign tm[1667] = 6423;
assign te[1667] = 14;
assign s[1668] = 2317652;
assign tm[1668] = 6421;
assign te[1668] = 14;
assign s[1669] = 2320860;
assign tm[1669] = 6419;
assign te[1669] = 14;
assign s[1670] = 2324068;
assign tm[1670] = 6417;
assign te[1670] = 14;
assign s[1671] = 2327275;
assign tm[1671] = 6415;
assign te[1671] = 14;
assign s[1672] = 2330481;
assign tm[1672] = 6413;
assign te[1672] = 14;
assign s[1673] = 2333686;
assign tm[1673] = 6411;
assign te[1673] = 14;
assign s[1674] = 2336890;
assign tm[1674] = 6409;
assign te[1674] = 14;
assign s[1675] = 2340093;
assign tm[1675] = 6408;
assign te[1675] = 14;
assign s[1676] = 2343295;
assign tm[1676] = 6406;
assign te[1676] = 14;
assign s[1677] = 2346497;
assign tm[1677] = 6404;
assign te[1677] = 14;
assign s[1678] = 2349696;
assign tm[1678] = 6402;
assign te[1678] = 14;
assign s[1679] = 2352896;
assign tm[1679] = 6400;
assign te[1679] = 14;
assign s[1680] = 2356094;
assign tm[1680] = 6398;
assign te[1680] = 14;
assign s[1681] = 2359291;
assign tm[1681] = 6396;
assign te[1681] = 14;
assign s[1682] = 2362488;
assign tm[1682] = 6394;
assign te[1682] = 14;
assign s[1683] = 2365684;
assign tm[1683] = 6392;
assign te[1683] = 14;
assign s[1684] = 2368878;
assign tm[1684] = 6390;
assign te[1684] = 14;
assign s[1685] = 2372072;
assign tm[1685] = 6389;
assign te[1685] = 14;
assign s[1686] = 2375264;
assign tm[1686] = 6387;
assign te[1686] = 14;
assign s[1687] = 2378456;
assign tm[1687] = 6385;
assign te[1687] = 14;
assign s[1688] = 2381647;
assign tm[1688] = 6383;
assign te[1688] = 14;
assign s[1689] = 2384836;
assign tm[1689] = 6381;
assign te[1689] = 14;
assign s[1690] = 2388025;
assign tm[1690] = 6379;
assign te[1690] = 14;
assign s[1691] = 2391213;
assign tm[1691] = 6377;
assign te[1691] = 14;
assign s[1692] = 2394400;
assign tm[1692] = 6375;
assign te[1692] = 14;
assign s[1693] = 2397586;
assign tm[1693] = 6373;
assign te[1693] = 14;
assign s[1694] = 2400771;
assign tm[1694] = 6371;
assign te[1694] = 14;
assign s[1695] = 2403955;
assign tm[1695] = 6370;
assign te[1695] = 14;
assign s[1696] = 2407139;
assign tm[1696] = 6368;
assign te[1696] = 14;
assign s[1697] = 2410320;
assign tm[1697] = 6366;
assign te[1697] = 14;
assign s[1698] = 2413502;
assign tm[1698] = 6364;
assign te[1698] = 14;
assign s[1699] = 2416683;
assign tm[1699] = 6362;
assign te[1699] = 14;
assign s[1700] = 2419862;
assign tm[1700] = 6360;
assign te[1700] = 14;
assign s[1701] = 2423040;
assign tm[1701] = 6358;
assign te[1701] = 14;
assign s[1702] = 2426218;
assign tm[1702] = 6356;
assign te[1702] = 14;
assign s[1703] = 2429395;
assign tm[1703] = 6355;
assign te[1703] = 14;
assign s[1704] = 2432570;
assign tm[1704] = 6353;
assign te[1704] = 14;
assign s[1705] = 2435745;
assign tm[1705] = 6351;
assign te[1705] = 14;
assign s[1706] = 2438919;
assign tm[1706] = 6349;
assign te[1706] = 14;
assign s[1707] = 2442091;
assign tm[1707] = 6347;
assign te[1707] = 14;
assign s[1708] = 2445264;
assign tm[1708] = 6345;
assign te[1708] = 14;
assign s[1709] = 2448434;
assign tm[1709] = 6343;
assign te[1709] = 14;
assign s[1710] = 2451604;
assign tm[1710] = 6342;
assign te[1710] = 14;
assign s[1711] = 2454774;
assign tm[1711] = 6340;
assign te[1711] = 14;
assign s[1712] = 2457942;
assign tm[1712] = 6338;
assign te[1712] = 14;
assign s[1713] = 2461109;
assign tm[1713] = 6336;
assign te[1713] = 14;
assign s[1714] = 2464276;
assign tm[1714] = 6334;
assign te[1714] = 14;
assign s[1715] = 2467441;
assign tm[1715] = 6332;
assign te[1715] = 14;
assign s[1716] = 2470606;
assign tm[1716] = 6330;
assign te[1716] = 14;
assign s[1717] = 2473770;
assign tm[1717] = 6329;
assign te[1717] = 14;
assign s[1718] = 2476932;
assign tm[1718] = 6327;
assign te[1718] = 14;
assign s[1719] = 2480094;
assign tm[1719] = 6325;
assign te[1719] = 14;
assign s[1720] = 2483255;
assign tm[1720] = 6323;
assign te[1720] = 14;
assign s[1721] = 2486415;
assign tm[1721] = 6321;
assign te[1721] = 14;
assign s[1722] = 2489574;
assign tm[1722] = 6319;
assign te[1722] = 14;
assign s[1723] = 2492732;
assign tm[1723] = 6318;
assign te[1723] = 14;
assign s[1724] = 2495889;
assign tm[1724] = 6316;
assign te[1724] = 14;
assign s[1725] = 2499046;
assign tm[1725] = 6314;
assign te[1725] = 14;
assign s[1726] = 2502201;
assign tm[1726] = 6312;
assign te[1726] = 14;
assign s[1727] = 2505356;
assign tm[1727] = 6310;
assign te[1727] = 14;
assign s[1728] = 2508510;
assign tm[1728] = 6308;
assign te[1728] = 14;
assign s[1729] = 2511661;
assign tm[1729] = 6307;
assign te[1729] = 14;
assign s[1730] = 2514814;
assign tm[1730] = 6305;
assign te[1730] = 14;
assign s[1731] = 2517964;
assign tm[1731] = 6303;
assign te[1731] = 14;
assign s[1732] = 2521114;
assign tm[1732] = 6301;
assign te[1732] = 14;
assign s[1733] = 2524263;
assign tm[1733] = 6299;
assign te[1733] = 14;
assign s[1734] = 2527411;
assign tm[1734] = 6298;
assign te[1734] = 14;
assign s[1735] = 2530558;
assign tm[1735] = 6296;
assign te[1735] = 14;
assign s[1736] = 2533705;
assign tm[1736] = 6294;
assign te[1736] = 14;
assign s[1737] = 2536851;
assign tm[1737] = 6292;
assign te[1737] = 14;
assign s[1738] = 2539994;
assign tm[1738] = 6290;
assign te[1738] = 14;
assign s[1739] = 2543138;
assign tm[1739] = 6288;
assign te[1739] = 14;
assign s[1740] = 2546281;
assign tm[1740] = 6287;
assign te[1740] = 14;
assign s[1741] = 2549423;
assign tm[1741] = 6285;
assign te[1741] = 14;
assign s[1742] = 2552564;
assign tm[1742] = 6283;
assign te[1742] = 14;
assign s[1743] = 2555704;
assign tm[1743] = 6281;
assign te[1743] = 14;
assign s[1744] = 2558842;
assign tm[1744] = 6279;
assign te[1744] = 14;
assign s[1745] = 2561981;
assign tm[1745] = 6278;
assign te[1745] = 14;
assign s[1746] = 2565118;
assign tm[1746] = 6276;
assign te[1746] = 14;
assign s[1747] = 2568255;
assign tm[1747] = 6274;
assign te[1747] = 14;
assign s[1748] = 2571389;
assign tm[1748] = 6272;
assign te[1748] = 14;
assign s[1749] = 2574525;
assign tm[1749] = 6270;
assign te[1749] = 14;
assign s[1750] = 2577658;
assign tm[1750] = 6269;
assign te[1750] = 14;
assign s[1751] = 2580791;
assign tm[1751] = 6267;
assign te[1751] = 14;
assign s[1752] = 2583923;
assign tm[1752] = 6265;
assign te[1752] = 14;
assign s[1753] = 2587053;
assign tm[1753] = 6263;
assign te[1753] = 14;
assign s[1754] = 2590184;
assign tm[1754] = 6261;
assign te[1754] = 14;
assign s[1755] = 2593313;
assign tm[1755] = 6260;
assign te[1755] = 14;
assign s[1756] = 2596441;
assign tm[1756] = 6258;
assign te[1756] = 14;
assign s[1757] = 2599568;
assign tm[1757] = 6256;
assign te[1757] = 14;
assign s[1758] = 2602695;
assign tm[1758] = 6254;
assign te[1758] = 14;
assign s[1759] = 2605820;
assign tm[1759] = 6253;
assign te[1759] = 14;
assign s[1760] = 2608946;
assign tm[1760] = 6251;
assign te[1760] = 14;
assign s[1761] = 2612069;
assign tm[1761] = 6249;
assign te[1761] = 14;
assign s[1762] = 2615193;
assign tm[1762] = 6247;
assign te[1762] = 14;
assign s[1763] = 2618314;
assign tm[1763] = 6245;
assign te[1763] = 14;
assign s[1764] = 2621436;
assign tm[1764] = 6244;
assign te[1764] = 14;
assign s[1765] = 2624556;
assign tm[1765] = 6242;
assign te[1765] = 14;
assign s[1766] = 2627676;
assign tm[1766] = 6240;
assign te[1766] = 14;
assign s[1767] = 2630794;
assign tm[1767] = 6238;
assign te[1767] = 14;
assign s[1768] = 2633912;
assign tm[1768] = 6237;
assign te[1768] = 14;
assign s[1769] = 2637029;
assign tm[1769] = 6235;
assign te[1769] = 14;
assign s[1770] = 2640144;
assign tm[1770] = 6233;
assign te[1770] = 14;
assign s[1771] = 2643259;
assign tm[1771] = 6231;
assign te[1771] = 14;
assign s[1772] = 2646374;
assign tm[1772] = 6230;
assign te[1772] = 14;
assign s[1773] = 2649486;
assign tm[1773] = 6228;
assign te[1773] = 14;
assign s[1774] = 2652600;
assign tm[1774] = 6226;
assign te[1774] = 14;
assign s[1775] = 2655711;
assign tm[1775] = 6224;
assign te[1775] = 14;
assign s[1776] = 2658821;
assign tm[1776] = 6223;
assign te[1776] = 14;
assign s[1777] = 2661932;
assign tm[1777] = 6221;
assign te[1777] = 14;
assign s[1778] = 2665040;
assign tm[1778] = 6219;
assign te[1778] = 14;
assign s[1779] = 2668148;
assign tm[1779] = 6217;
assign te[1779] = 14;
assign s[1780] = 2671255;
assign tm[1780] = 6216;
assign te[1780] = 14;
assign s[1781] = 2674361;
assign tm[1781] = 6214;
assign te[1781] = 14;
assign s[1782] = 2677467;
assign tm[1782] = 6212;
assign te[1782] = 14;
assign s[1783] = 2680571;
assign tm[1783] = 6210;
assign te[1783] = 14;
assign s[1784] = 2683675;
assign tm[1784] = 6209;
assign te[1784] = 14;
assign s[1785] = 2686778;
assign tm[1785] = 6207;
assign te[1785] = 14;
assign s[1786] = 2689880;
assign tm[1786] = 6205;
assign te[1786] = 14;
assign s[1787] = 2692981;
assign tm[1787] = 6203;
assign te[1787] = 14;
assign s[1788] = 2696081;
assign tm[1788] = 6202;
assign te[1788] = 14;
assign s[1789] = 2699180;
assign tm[1789] = 6200;
assign te[1789] = 14;
assign s[1790] = 2702279;
assign tm[1790] = 6198;
assign te[1790] = 14;
assign s[1791] = 2705377;
assign tm[1791] = 6196;
assign te[1791] = 14;
assign s[1792] = 2708473;
assign tm[1792] = 6195;
assign te[1792] = 14;
assign s[1793] = 2711569;
assign tm[1793] = 6193;
assign te[1793] = 14;
assign s[1794] = 2714663;
assign tm[1794] = 6191;
assign te[1794] = 14;
assign s[1795] = 2717758;
assign tm[1795] = 6189;
assign te[1795] = 14;
assign s[1796] = 2720851;
assign tm[1796] = 6188;
assign te[1796] = 14;
assign s[1797] = 2723944;
assign tm[1797] = 6186;
assign te[1797] = 14;
assign s[1798] = 2727035;
assign tm[1798] = 6184;
assign te[1798] = 14;
assign s[1799] = 2730126;
assign tm[1799] = 6183;
assign te[1799] = 14;
assign s[1800] = 2733215;
assign tm[1800] = 6181;
assign te[1800] = 14;
assign s[1801] = 2736305;
assign tm[1801] = 6179;
assign te[1801] = 14;
assign s[1802] = 2739392;
assign tm[1802] = 6177;
assign te[1802] = 14;
assign s[1803] = 2742480;
assign tm[1803] = 6176;
assign te[1803] = 14;
assign s[1804] = 2745567;
assign tm[1804] = 6174;
assign te[1804] = 14;
assign s[1805] = 2748652;
assign tm[1805] = 6172;
assign te[1805] = 14;
assign s[1806] = 2751737;
assign tm[1806] = 6171;
assign te[1806] = 14;
assign s[1807] = 2754820;
assign tm[1807] = 6169;
assign te[1807] = 14;
assign s[1808] = 2757903;
assign tm[1808] = 6167;
assign te[1808] = 14;
assign s[1809] = 2760986;
assign tm[1809] = 6165;
assign te[1809] = 14;
assign s[1810] = 2764067;
assign tm[1810] = 6164;
assign te[1810] = 14;
assign s[1811] = 2767147;
assign tm[1811] = 6162;
assign te[1811] = 14;
assign s[1812] = 2770227;
assign tm[1812] = 6160;
assign te[1812] = 14;
assign s[1813] = 2773306;
assign tm[1813] = 6159;
assign te[1813] = 14;
assign s[1814] = 2776383;
assign tm[1814] = 6157;
assign te[1814] = 14;
assign s[1815] = 2779460;
assign tm[1815] = 6155;
assign te[1815] = 14;
assign s[1816] = 2782537;
assign tm[1816] = 6154;
assign te[1816] = 14;
assign s[1817] = 2785612;
assign tm[1817] = 6152;
assign te[1817] = 14;
assign s[1818] = 2788686;
assign tm[1818] = 6150;
assign te[1818] = 14;
assign s[1819] = 2791760;
assign tm[1819] = 6148;
assign te[1819] = 14;
assign s[1820] = 2794833;
assign tm[1820] = 6147;
assign te[1820] = 14;
assign s[1821] = 2797905;
assign tm[1821] = 6145;
assign te[1821] = 14;
assign s[1822] = 2800976;
assign tm[1822] = 6143;
assign te[1822] = 14;
assign s[1823] = 2804046;
assign tm[1823] = 6142;
assign te[1823] = 14;
assign s[1824] = 2807116;
assign tm[1824] = 6140;
assign te[1824] = 14;
assign s[1825] = 2810184;
assign tm[1825] = 6138;
assign te[1825] = 14;
assign s[1826] = 2813252;
assign tm[1826] = 6137;
assign te[1826] = 14;
assign s[1827] = 2816319;
assign tm[1827] = 6135;
assign te[1827] = 14;
assign s[1828] = 2819385;
assign tm[1828] = 6133;
assign te[1828] = 14;
assign s[1829] = 2822450;
assign tm[1829] = 6132;
assign te[1829] = 14;
assign s[1830] = 2825514;
assign tm[1830] = 6130;
assign te[1830] = 14;
assign s[1831] = 2828578;
assign tm[1831] = 6128;
assign te[1831] = 14;
assign s[1832] = 2831641;
assign tm[1832] = 6127;
assign te[1832] = 14;
assign s[1833] = 2834703;
assign tm[1833] = 6125;
assign te[1833] = 14;
assign s[1834] = 2837763;
assign tm[1834] = 6123;
assign te[1834] = 14;
assign s[1835] = 2840824;
assign tm[1835] = 6122;
assign te[1835] = 14;
assign s[1836] = 2843884;
assign tm[1836] = 6120;
assign te[1836] = 14;
assign s[1837] = 2846942;
assign tm[1837] = 6118;
assign te[1837] = 14;
assign s[1838] = 2849999;
assign tm[1838] = 6117;
assign te[1838] = 14;
assign s[1839] = 2853056;
assign tm[1839] = 6115;
assign te[1839] = 14;
assign s[1840] = 2856113;
assign tm[1840] = 6113;
assign te[1840] = 14;
assign s[1841] = 2859168;
assign tm[1841] = 6112;
assign te[1841] = 14;
assign s[1842] = 2862223;
assign tm[1842] = 6110;
assign te[1842] = 14;
assign s[1843] = 2865276;
assign tm[1843] = 6108;
assign te[1843] = 14;
assign s[1844] = 2868328;
assign tm[1844] = 6107;
assign te[1844] = 14;
assign s[1845] = 2871380;
assign tm[1845] = 6105;
assign te[1845] = 14;
assign s[1846] = 2874431;
assign tm[1846] = 6103;
assign te[1846] = 14;
assign s[1847] = 2877482;
assign tm[1847] = 6102;
assign te[1847] = 14;
assign s[1848] = 2880531;
assign tm[1848] = 6100;
assign te[1848] = 14;
assign s[1849] = 2883579;
assign tm[1849] = 6098;
assign te[1849] = 14;
assign s[1850] = 2886627;
assign tm[1850] = 6097;
assign te[1850] = 14;
assign s[1851] = 2889675;
assign tm[1851] = 6095;
assign te[1851] = 14;
assign s[1852] = 2892720;
assign tm[1852] = 6093;
assign te[1852] = 14;
assign s[1853] = 2895766;
assign tm[1853] = 6092;
assign te[1853] = 14;
assign s[1854] = 2898810;
assign tm[1854] = 6090;
assign te[1854] = 14;
assign s[1855] = 2901854;
assign tm[1855] = 6088;
assign te[1855] = 14;
assign s[1856] = 2904897;
assign tm[1856] = 6087;
assign te[1856] = 14;
assign s[1857] = 2907939;
assign tm[1857] = 6085;
assign te[1857] = 14;
assign s[1858] = 2910980;
assign tm[1858] = 6084;
assign te[1858] = 14;
assign s[1859] = 2914021;
assign tm[1859] = 6082;
assign te[1859] = 14;
assign s[1860] = 2917060;
assign tm[1860] = 6080;
assign te[1860] = 14;
assign s[1861] = 2920099;
assign tm[1861] = 6079;
assign te[1861] = 14;
assign s[1862] = 2923137;
assign tm[1862] = 6077;
assign te[1862] = 14;
assign s[1863] = 2926174;
assign tm[1863] = 6075;
assign te[1863] = 14;
assign s[1864] = 2929210;
assign tm[1864] = 6074;
assign te[1864] = 14;
assign s[1865] = 2932246;
assign tm[1865] = 6072;
assign te[1865] = 14;
assign s[1866] = 2935280;
assign tm[1866] = 6070;
assign te[1866] = 14;
assign s[1867] = 2938314;
assign tm[1867] = 6069;
assign te[1867] = 14;
assign s[1868] = 2941348;
assign tm[1868] = 6067;
assign te[1868] = 14;
assign s[1869] = 2944379;
assign tm[1869] = 6066;
assign te[1869] = 14;
assign s[1870] = 2947410;
assign tm[1870] = 6064;
assign te[1870] = 14;
assign s[1871] = 2950441;
assign tm[1871] = 6062;
assign te[1871] = 14;
assign s[1872] = 2953471;
assign tm[1872] = 6061;
assign te[1872] = 14;
assign s[1873] = 2956500;
assign tm[1873] = 6059;
assign te[1873] = 14;
assign s[1874] = 2959528;
assign tm[1874] = 6057;
assign te[1874] = 14;
assign s[1875] = 2962556;
assign tm[1875] = 6056;
assign te[1875] = 14;
assign s[1876] = 2965583;
assign tm[1876] = 6054;
assign te[1876] = 14;
assign s[1877] = 2968608;
assign tm[1877] = 6053;
assign te[1877] = 14;
assign s[1878] = 2971634;
assign tm[1878] = 6051;
assign te[1878] = 14;
assign s[1879] = 2974657;
assign tm[1879] = 6049;
assign te[1879] = 14;
assign s[1880] = 2977681;
assign tm[1880] = 6048;
assign te[1880] = 14;
assign s[1881] = 2980703;
assign tm[1881] = 6046;
assign te[1881] = 14;
assign s[1882] = 2983725;
assign tm[1882] = 6045;
assign te[1882] = 14;
assign s[1883] = 2986746;
assign tm[1883] = 6043;
assign te[1883] = 14;
assign s[1884] = 2989766;
assign tm[1884] = 6041;
assign te[1884] = 14;
assign s[1885] = 2992785;
assign tm[1885] = 6040;
assign te[1885] = 14;
assign s[1886] = 2995804;
assign tm[1886] = 6038;
assign te[1886] = 14;
assign s[1887] = 2998822;
assign tm[1887] = 6037;
assign te[1887] = 14;
assign s[1888] = 3001838;
assign tm[1888] = 6035;
assign te[1888] = 14;
assign s[1889] = 3004855;
assign tm[1889] = 6033;
assign te[1889] = 14;
assign s[1890] = 3007870;
assign tm[1890] = 6032;
assign te[1890] = 14;
assign s[1891] = 3010884;
assign tm[1891] = 6030;
assign te[1891] = 14;
assign s[1892] = 3013898;
assign tm[1892] = 6029;
assign te[1892] = 14;
assign s[1893] = 3016912;
assign tm[1893] = 6027;
assign te[1893] = 14;
assign s[1894] = 3019923;
assign tm[1894] = 6025;
assign te[1894] = 14;
assign s[1895] = 3022935;
assign tm[1895] = 6024;
assign te[1895] = 14;
assign s[1896] = 3025945;
assign tm[1896] = 6022;
assign te[1896] = 14;
assign s[1897] = 3028955;
assign tm[1897] = 6021;
assign te[1897] = 14;
assign s[1898] = 3031965;
assign tm[1898] = 6019;
assign te[1898] = 14;
assign s[1899] = 3034972;
assign tm[1899] = 6017;
assign te[1899] = 14;
assign s[1900] = 3037980;
assign tm[1900] = 6016;
assign te[1900] = 14;
assign s[1901] = 3040986;
assign tm[1901] = 6014;
assign te[1901] = 14;
assign s[1902] = 3043992;
assign tm[1902] = 6013;
assign te[1902] = 14;
assign s[1903] = 3046998;
assign tm[1903] = 6011;
assign te[1903] = 14;
assign s[1904] = 3050001;
assign tm[1904] = 6010;
assign te[1904] = 14;
assign s[1905] = 3053005;
assign tm[1905] = 6008;
assign te[1905] = 14;
assign s[1906] = 3056008;
assign tm[1906] = 6006;
assign te[1906] = 14;
assign s[1907] = 3059009;
assign tm[1907] = 6005;
assign te[1907] = 14;
assign s[1908] = 3062010;
assign tm[1908] = 6003;
assign te[1908] = 14;
assign s[1909] = 3065010;
assign tm[1909] = 6002;
assign te[1909] = 14;
assign s[1910] = 3068010;
assign tm[1910] = 6000;
assign te[1910] = 14;
assign s[1911] = 3071009;
assign tm[1911] = 5999;
assign te[1911] = 14;
assign s[1912] = 3074007;
assign tm[1912] = 5997;
assign te[1912] = 14;
assign s[1913] = 3077004;
assign tm[1913] = 5995;
assign te[1913] = 14;
assign s[1914] = 3080000;
assign tm[1914] = 5994;
assign te[1914] = 14;
assign s[1915] = 3082996;
assign tm[1915] = 5992;
assign te[1915] = 14;
assign s[1916] = 3085990;
assign tm[1916] = 5991;
assign te[1916] = 14;
assign s[1917] = 3088985;
assign tm[1917] = 5989;
assign te[1917] = 14;
assign s[1918] = 3091978;
assign tm[1918] = 5988;
assign te[1918] = 14;
assign s[1919] = 3094971;
assign tm[1919] = 5986;
assign te[1919] = 14;
assign s[1920] = 3097962;
assign tm[1920] = 5984;
assign te[1920] = 14;
assign s[1921] = 3100953;
assign tm[1921] = 5983;
assign te[1921] = 14;
assign s[1922] = 3103943;
assign tm[1922] = 5981;
assign te[1922] = 14;
assign s[1923] = 3106933;
assign tm[1923] = 5980;
assign te[1923] = 14;
assign s[1924] = 3109921;
assign tm[1924] = 5978;
assign te[1924] = 14;
assign s[1925] = 3112909;
assign tm[1925] = 5977;
assign te[1925] = 14;
assign s[1926] = 3115897;
assign tm[1926] = 5975;
assign te[1926] = 14;
assign s[1927] = 3118882;
assign tm[1927] = 5974;
assign te[1927] = 14;
assign s[1928] = 3121868;
assign tm[1928] = 5972;
assign te[1928] = 14;
assign s[1929] = 3124852;
assign tm[1929] = 5970;
assign te[1929] = 14;
assign s[1930] = 3127837;
assign tm[1930] = 5969;
assign te[1930] = 14;
assign s[1931] = 3130820;
assign tm[1931] = 5967;
assign te[1931] = 14;
assign s[1932] = 3133802;
assign tm[1932] = 5966;
assign te[1932] = 14;
assign s[1933] = 3136784;
assign tm[1933] = 5964;
assign te[1933] = 14;
assign s[1934] = 3139764;
assign tm[1934] = 5963;
assign te[1934] = 14;
assign s[1935] = 3142745;
assign tm[1935] = 5961;
assign te[1935] = 14;
assign s[1936] = 3145723;
assign tm[1936] = 5960;
assign te[1936] = 14;
assign s[1937] = 3148702;
assign tm[1937] = 5958;
assign te[1937] = 14;
assign s[1938] = 3151680;
assign tm[1938] = 5957;
assign te[1938] = 14;
assign s[1939] = 3154657;
assign tm[1939] = 5955;
assign te[1939] = 14;
assign s[1940] = 3157633;
assign tm[1940] = 5953;
assign te[1940] = 14;
assign s[1941] = 3160609;
assign tm[1941] = 5952;
assign te[1941] = 14;
assign s[1942] = 3163583;
assign tm[1942] = 5950;
assign te[1942] = 14;
assign s[1943] = 3166557;
assign tm[1943] = 5949;
assign te[1943] = 14;
assign s[1944] = 3169530;
assign tm[1944] = 5947;
assign te[1944] = 14;
assign s[1945] = 3172503;
assign tm[1945] = 5946;
assign te[1945] = 14;
assign s[1946] = 3175474;
assign tm[1946] = 5944;
assign te[1946] = 14;
assign s[1947] = 3178445;
assign tm[1947] = 5943;
assign te[1947] = 14;
assign s[1948] = 3181415;
assign tm[1948] = 5941;
assign te[1948] = 14;
assign s[1949] = 3184385;
assign tm[1949] = 5940;
assign te[1949] = 14;
assign s[1950] = 3187354;
assign tm[1950] = 5938;
assign te[1950] = 14;
assign s[1951] = 3190321;
assign tm[1951] = 5937;
assign te[1951] = 14;
assign s[1952] = 3193288;
assign tm[1952] = 5935;
assign te[1952] = 14;
assign s[1953] = 3196255;
assign tm[1953] = 5934;
assign te[1953] = 14;
assign s[1954] = 3199220;
assign tm[1954] = 5932;
assign te[1954] = 14;
assign s[1955] = 3202185;
assign tm[1955] = 5931;
assign te[1955] = 14;
assign s[1956] = 3205149;
assign tm[1956] = 5929;
assign te[1956] = 14;
assign s[1957] = 3208112;
assign tm[1957] = 5928;
assign te[1957] = 14;
assign s[1958] = 3211074;
assign tm[1958] = 5926;
assign te[1958] = 14;
assign s[1959] = 3214037;
assign tm[1959] = 5925;
assign te[1959] = 14;
assign s[1960] = 3216998;
assign tm[1960] = 5923;
assign te[1960] = 14;
assign s[1961] = 3219958;
assign tm[1961] = 5921;
assign te[1961] = 14;
assign s[1962] = 3222917;
assign tm[1962] = 5920;
assign te[1962] = 14;
assign s[1963] = 3225876;
assign tm[1963] = 5918;
assign te[1963] = 14;
assign s[1964] = 3228834;
assign tm[1964] = 5917;
assign te[1964] = 14;
assign s[1965] = 3231791;
assign tm[1965] = 5915;
assign te[1965] = 14;
assign s[1966] = 3234747;
assign tm[1966] = 5914;
assign te[1966] = 14;
assign s[1967] = 3237704;
assign tm[1967] = 5912;
assign te[1967] = 14;
assign s[1968] = 3240658;
assign tm[1968] = 5911;
assign te[1968] = 14;
assign s[1969] = 3243613;
assign tm[1969] = 5909;
assign te[1969] = 14;
assign s[1970] = 3246565;
assign tm[1970] = 5908;
assign te[1970] = 14;
assign s[1971] = 3249519;
assign tm[1971] = 5906;
assign te[1971] = 14;
assign s[1972] = 3252471;
assign tm[1972] = 5905;
assign te[1972] = 14;
assign s[1973] = 3255422;
assign tm[1973] = 5903;
assign te[1973] = 14;
assign s[1974] = 3258372;
assign tm[1974] = 5902;
assign te[1974] = 14;
assign s[1975] = 3261322;
assign tm[1975] = 5900;
assign te[1975] = 14;
assign s[1976] = 3264271;
assign tm[1976] = 5899;
assign te[1976] = 14;
assign s[1977] = 3267219;
assign tm[1977] = 5897;
assign te[1977] = 14;
assign s[1978] = 3270166;
assign tm[1978] = 5896;
assign te[1978] = 14;
assign s[1979] = 3273113;
assign tm[1979] = 5894;
assign te[1979] = 14;
assign s[1980] = 3276059;
assign tm[1980] = 5893;
assign te[1980] = 14;
assign s[1981] = 3279005;
assign tm[1981] = 5891;
assign te[1981] = 14;
assign s[1982] = 3281949;
assign tm[1982] = 5890;
assign te[1982] = 14;
assign s[1983] = 3284893;
assign tm[1983] = 5889;
assign te[1983] = 14;
assign s[1984] = 3287836;
assign tm[1984] = 5887;
assign te[1984] = 14;
assign s[1985] = 3290779;
assign tm[1985] = 5886;
assign te[1985] = 14;
assign s[1986] = 3293720;
assign tm[1986] = 5884;
assign te[1986] = 14;
assign s[1987] = 3296660;
assign tm[1987] = 5883;
assign te[1987] = 14;
assign s[1988] = 3299601;
assign tm[1988] = 5881;
assign te[1988] = 14;
assign s[1989] = 3302540;
assign tm[1989] = 5880;
assign te[1989] = 14;
assign s[1990] = 3305478;
assign tm[1990] = 5878;
assign te[1990] = 14;
assign s[1991] = 3308416;
assign tm[1991] = 5877;
assign te[1991] = 14;
assign s[1992] = 3311353;
assign tm[1992] = 5875;
assign te[1992] = 14;
assign s[1993] = 3314290;
assign tm[1993] = 5874;
assign te[1993] = 14;
assign s[1994] = 3317225;
assign tm[1994] = 5872;
assign te[1994] = 14;
assign s[1995] = 3320160;
assign tm[1995] = 5871;
assign te[1995] = 14;
assign s[1996] = 3323094;
assign tm[1996] = 5869;
assign te[1996] = 14;
assign s[1997] = 3326028;
assign tm[1997] = 5868;
assign te[1997] = 14;
assign s[1998] = 3328961;
assign tm[1998] = 5866;
assign te[1998] = 14;
assign s[1999] = 3331892;
assign tm[1999] = 5865;
assign te[1999] = 14;
assign s[2000] = 3334824;
assign tm[2000] = 5863;
assign te[2000] = 14;
assign s[2001] = 3337754;
assign tm[2001] = 5862;
assign te[2001] = 14;
assign s[2002] = 3340684;
assign tm[2002] = 5860;
assign te[2002] = 14;
assign s[2003] = 3343613;
assign tm[2003] = 5859;
assign te[2003] = 14;
assign s[2004] = 3346542;
assign tm[2004] = 5858;
assign te[2004] = 14;
assign s[2005] = 3349469;
assign tm[2005] = 5856;
assign te[2005] = 14;
assign s[2006] = 3352396;
assign tm[2006] = 5855;
assign te[2006] = 14;
assign s[2007] = 3355322;
assign tm[2007] = 5853;
assign te[2007] = 14;
assign s[2008] = 3358247;
assign tm[2008] = 5852;
assign te[2008] = 14;
assign s[2009] = 3361172;
assign tm[2009] = 5850;
assign te[2009] = 14;
assign s[2010] = 3364096;
assign tm[2010] = 5849;
assign te[2010] = 14;
assign s[2011] = 3367019;
assign tm[2011] = 5847;
assign te[2011] = 14;
assign s[2012] = 3369941;
assign tm[2012] = 5846;
assign te[2012] = 14;
assign s[2013] = 3372863;
assign tm[2013] = 5844;
assign te[2013] = 14;
assign s[2014] = 3375785;
assign tm[2014] = 5843;
assign te[2014] = 14;
assign s[2015] = 3378705;
assign tm[2015] = 5842;
assign te[2015] = 14;
assign s[2016] = 3381625;
assign tm[2016] = 5840;
assign te[2016] = 14;
assign s[2017] = 3384543;
assign tm[2017] = 5839;
assign te[2017] = 14;
assign s[2018] = 3387461;
assign tm[2018] = 5837;
assign te[2018] = 14;
assign s[2019] = 3390378;
assign tm[2019] = 5836;
assign te[2019] = 14;
assign s[2020] = 3393295;
assign tm[2020] = 5834;
assign te[2020] = 14;
assign s[2021] = 3396212;
assign tm[2021] = 5833;
assign te[2021] = 14;
assign s[2022] = 3399126;
assign tm[2022] = 5831;
assign te[2022] = 14;
assign s[2023] = 3402041;
assign tm[2023] = 5830;
assign te[2023] = 14;
assign s[2024] = 3404955;
assign tm[2024] = 5829;
assign te[2024] = 14;
assign s[2025] = 3407867;
assign tm[2025] = 5827;
assign te[2025] = 14;
assign s[2026] = 3410780;
assign tm[2026] = 5826;
assign te[2026] = 14;
assign s[2027] = 3413692;
assign tm[2027] = 5824;
assign te[2027] = 14;
assign s[2028] = 3416603;
assign tm[2028] = 5823;
assign te[2028] = 14;
assign s[2029] = 3419513;
assign tm[2029] = 5821;
assign te[2029] = 14;
assign s[2030] = 3422423;
assign tm[2030] = 5820;
assign te[2030] = 14;
assign s[2031] = 3425331;
assign tm[2031] = 5818;
assign te[2031] = 14;
assign s[2032] = 3428239;
assign tm[2032] = 5817;
assign te[2032] = 14;
assign s[2033] = 3431147;
assign tm[2033] = 5816;
assign te[2033] = 14;
assign s[2034] = 3434053;
assign tm[2034] = 5814;
assign te[2034] = 14;
assign s[2035] = 3436959;
assign tm[2035] = 5813;
assign te[2035] = 14;
assign s[2036] = 3439864;
assign tm[2036] = 5811;
assign te[2036] = 14;
assign s[2037] = 3442768;
assign tm[2037] = 5810;
assign te[2037] = 14;
assign s[2038] = 3445672;
assign tm[2038] = 5808;
assign te[2038] = 14;
assign s[2039] = 3448576;
assign tm[2039] = 5807;
assign te[2039] = 14;
assign s[2040] = 3451478;
assign tm[2040] = 5806;
assign te[2040] = 14;
assign s[2041] = 3454379;
assign tm[2041] = 5804;
assign te[2041] = 14;
assign s[2042] = 3457280;
assign tm[2042] = 5803;
assign te[2042] = 14;
assign s[2043] = 3460181;
assign tm[2043] = 5801;
assign te[2043] = 14;
assign s[2044] = 3463081;
assign tm[2044] = 5800;
assign te[2044] = 14;
assign s[2045] = 3465979;
assign tm[2045] = 5798;
assign te[2045] = 14;
assign s[2046] = 3468877;
assign tm[2046] = 5797;
assign te[2046] = 14;
assign s[2047] = 3471775;
assign tm[2047] = 5796;
assign te[2047] = 14;

wire [8:0] se;
assign se = adata[23] ? {1'b0,((adata[30:23] >> 1) + 8'd64)} : {1'b0,((adata[30:23] >> 1) + 8'd63)};

wire [10:0] key;
assign key = adata[23:13];

wire [25:0] ta;
assign ta = tm[key] * adata[12:0];

reg [25:0] ta_reg;
(* ram_style = "distributed" *) reg [5:0] te_reg;
(* ram_style = "distributed" *) reg [22:0] s_reg;
reg notzero_reg;
reg [8:0] se_reg;
reg flag_reg;
reg [4:0] address_reg;
always_ff@(posedge clk) begin
ta_reg <= ta;
te_reg <= te[key];
s_reg <= s[key];
notzero_reg <= |adata[30:23];
se_reg <= se;
flag_reg <= flag_in;
address_reg <= address_in;
end

wire [12:0] ta_s;
assign ta_s = ta_reg >> te_reg;

wire [22:0] kari;
assign kari = s_reg + ta_s;

always_ff@(posedge clk) begin
result <= notzero_reg ? {se_reg,kari} : 0;
flag_out <= flag_reg;
address_out <= address_reg;
end  

endmodule

`default_nettype wire
