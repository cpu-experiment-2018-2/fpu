`default_nettype none

module fsqrt(
input wire [31:0] adata,
output reg [31:0] result,
input wire clk,
input wire flag_in,
input wire [4:0] address_in,
output reg flag_out,
output reg [4:0] address_out);

(* ram_style = "distributed" *) reg [22:0] key [511:0];
(* ram_style = "distributed" *) reg [13:0] key2 [511:0];

assign key[0] = 3474675;
assign key2[0] = 11585;
assign key[1] = 3497823;
assign key2[1] = 11562;
assign key[2] = 3520926;
assign key2[2] = 11540;
assign key[3] = 3543984;
assign key2[3] = 11517;
assign key[4] = 3566998;
assign key2[4] = 11495;
assign key[5] = 3589967;
assign key2[5] = 11473;
assign key[6] = 3612893;
assign key2[6] = 11451;
assign key[7] = 3635775;
assign key2[7] = 11430;
assign key[8] = 3658613;
assign key2[8] = 11408;
assign key[9] = 3681408;
assign key2[9] = 11386;
assign key[10] = 3704160;
assign key2[10] = 11365;
assign key[11] = 3726870;
assign key2[11] = 11344;
assign key[12] = 3749537;
assign key2[12] = 11322;
assign key[13] = 3772161;
assign key2[13] = 11301;
assign key[14] = 3794744;
assign key2[14] = 11280;
assign key[15] = 3817285;
assign key2[15] = 11260;
assign key[16] = 3839784;
assign key2[16] = 11239;
assign key[17] = 3862242;
assign key2[17] = 11218;
assign key[18] = 3884659;
assign key2[18] = 11198;
assign key[19] = 3907035;
assign key2[19] = 11177;
assign key[20] = 3929371;
assign key2[20] = 11157;
assign key[21] = 3951666;
assign key2[21] = 11137;
assign key[22] = 3973921;
assign key2[22] = 11117;
assign key[23] = 3996136;
assign key2[23] = 11097;
assign key[24] = 4018311;
assign key2[24] = 11077;
assign key[25] = 4040446;
assign key2[25] = 11057;
assign key[26] = 4062542;
assign key2[26] = 11038;
assign key[27] = 4084599;
assign key2[27] = 11018;
assign key[28] = 4106617;
assign key2[28] = 10999;
assign key[29] = 4128596;
assign key2[29] = 10980;
assign key[30] = 4150537;
assign key2[30] = 10960;
assign key[31] = 4172440;
assign key2[31] = 10941;
assign key[32] = 4194304;
assign key2[32] = 10922;
assign key[33] = 4216130;
assign key2[33] = 10903;
assign key[34] = 4237919;
assign key2[34] = 10884;
assign key[35] = 4259670;
assign key2[35] = 10866;
assign key[36] = 4281384;
assign key2[36] = 10847;
assign key[37] = 4303061;
assign key2[37] = 10829;
assign key[38] = 4324700;
assign key2[38] = 10810;
assign key[39] = 4346303;
assign key2[39] = 10792;
assign key[40] = 4367870;
assign key2[40] = 10774;
assign key[41] = 4389400;
assign key2[41] = 10755;
assign key[42] = 4410893;
assign key2[42] = 10737;
assign key[43] = 4432351;
assign key2[43] = 10719;
assign key[44] = 4453773;
assign key2[44] = 10701;
assign key[45] = 4475159;
assign key2[45] = 10684;
assign key[46] = 4496510;
assign key2[46] = 10666;
assign key[47] = 4517825;
assign key2[47] = 10648;
assign key[48] = 4539105;
assign key2[48] = 10631;
assign key[49] = 4560350;
assign key2[49] = 10613;
assign key[50] = 4581561;
assign key2[50] = 10596;
assign key[51] = 4602737;
assign key2[51] = 10579;
assign key[52] = 4623878;
assign key2[52] = 10562;
assign key[53] = 4644985;
assign key2[53] = 10544;
assign key[54] = 4666058;
assign key2[54] = 10527;
assign key[55] = 4687097;
assign key2[55] = 10511;
assign key[56] = 4708102;
assign key2[56] = 10494;
assign key[57] = 4729074;
assign key2[57] = 10477;
assign key[58] = 4750012;
assign key2[58] = 10460;
assign key[59] = 4770916;
assign key2[59] = 10444;
assign key[60] = 4791788;
assign key2[60] = 10427;
assign key[61] = 4812627;
assign key2[61] = 10411;
assign key[62] = 4833432;
assign key2[62] = 10394;
assign key[63] = 4854205;
assign key2[63] = 10378;
assign key[64] = 4874946;
assign key2[64] = 10362;
assign key[65] = 4895654;
assign key2[65] = 10345;
assign key[66] = 4916330;
assign key2[66] = 10329;
assign key[67] = 4936974;
assign key2[67] = 10313;
assign key[68] = 4957586;
assign key2[68] = 10297;
assign key[69] = 4978166;
assign key2[69] = 10282;
assign key[70] = 4998714;
assign key2[70] = 10266;
assign key[71] = 5019231;
assign key2[71] = 10250;
assign key[72] = 5039717;
assign key2[72] = 10235;
assign key[73] = 5060171;
assign key2[73] = 10219;
assign key[74] = 5080595;
assign key2[74] = 10203;
assign key[75] = 5100987;
assign key2[75] = 10188;
assign key[76] = 5121349;
assign key2[76] = 10173;
assign key[77] = 5141680;
assign key2[77] = 10157;
assign key[78] = 5161980;
assign key2[78] = 10142;
assign key[79] = 5182250;
assign key2[79] = 10127;
assign key[80] = 5202490;
assign key2[80] = 10112;
assign key[81] = 5222700;
assign key2[81] = 10097;
assign key[82] = 5242880;
assign key2[82] = 10082;
assign key[83] = 5263030;
assign key2[83] = 10067;
assign key[84] = 5283150;
assign key2[84] = 10052;
assign key[85] = 5303241;
assign key2[85] = 10038;
assign key[86] = 5323302;
assign key2[86] = 10023;
assign key[87] = 5343334;
assign key2[87] = 10008;
assign key[88] = 5363337;
assign key2[88] = 9994;
assign key[89] = 5383311;
assign key2[89] = 9979;
assign key[90] = 5403256;
assign key2[90] = 9965;
assign key[91] = 5423172;
assign key2[91] = 9950;
assign key[92] = 5443059;
assign key2[92] = 9936;
assign key[93] = 5462918;
assign key2[93] = 9922;
assign key[94] = 5482749;
assign key2[94] = 9908;
assign key[95] = 5502551;
assign key2[95] = 9893;
assign key[96] = 5522325;
assign key2[96] = 9879;
assign key[97] = 5542070;
assign key2[97] = 9865;
assign key[98] = 5561788;
assign key2[98] = 9851;
assign key[99] = 5581478;
assign key2[99] = 9838;
assign key[100] = 5601141;
assign key2[100] = 9824;
assign key[101] = 5620775;
assign key2[101] = 9810;
assign key[102] = 5640383;
assign key2[102] = 9796;
assign key[103] = 5659963;
assign key2[103] = 9783;
assign key[104] = 5679515;
assign key2[104] = 9769;
assign key[105] = 5699041;
assign key2[105] = 9755;
assign key[106] = 5718539;
assign key2[106] = 9742;
assign key[107] = 5738011;
assign key2[107] = 9729;
assign key[108] = 5757456;
assign key2[108] = 9715;
assign key[109] = 5776874;
assign key2[109] = 9702;
assign key[110] = 5796265;
assign key2[110] = 9689;
assign key[111] = 5815630;
assign key2[111] = 9675;
assign key[112] = 5834969;
assign key2[112] = 9662;
assign key[113] = 5854281;
assign key2[113] = 9649;
assign key[114] = 5873568;
assign key2[114] = 9636;
assign key[115] = 5892828;
assign key2[115] = 9623;
assign key[116] = 5912062;
assign key2[116] = 9610;
assign key[117] = 5931270;
assign key2[117] = 9597;
assign key[118] = 5950453;
assign key2[118] = 9584;
assign key[119] = 5969610;
assign key2[119] = 9572;
assign key[120] = 5988742;
assign key2[120] = 9559;
assign key[121] = 6007848;
assign key2[121] = 9546;
assign key[122] = 6026929;
assign key2[122] = 9534;
assign key[123] = 6045984;
assign key2[123] = 9521;
assign key[124] = 6065015;
assign key2[124] = 9508;
assign key[125] = 6084020;
assign key2[125] = 9496;
assign key[126] = 6103001;
assign key2[126] = 9484;
assign key[127] = 6121956;
assign key2[127] = 9471;
assign key[128] = 6140887;
assign key2[128] = 9459;
assign key[129] = 6159794;
assign key2[129] = 9447;
assign key[130] = 6178675;
assign key2[130] = 9434;
assign key[131] = 6197533;
assign key2[131] = 9422;
assign key[132] = 6216366;
assign key2[132] = 9410;
assign key[133] = 6235174;
assign key2[133] = 9398;
assign key[134] = 6253959;
assign key2[134] = 9386;
assign key[135] = 6272719;
assign key2[135] = 9374;
assign key[136] = 6291456;
assign key2[136] = 9362;
assign key[137] = 6310169;
assign key2[137] = 9350;
assign key[138] = 6328857;
assign key2[138] = 9338;
assign key[139] = 6347523;
assign key2[139] = 9326;
assign key[140] = 6366164;
assign key2[140] = 9314;
assign key[141] = 6384782;
assign key2[141] = 9303;
assign key[142] = 6403377;
assign key2[142] = 9291;
assign key[143] = 6421948;
assign key2[143] = 9279;
assign key[144] = 6440496;
assign key2[144] = 9268;
assign key[145] = 6459021;
assign key2[145] = 9256;
assign key[146] = 6477523;
assign key2[146] = 9245;
assign key[147] = 6496001;
assign key2[147] = 9233;
assign key[148] = 6514457;
assign key2[148] = 9222;
assign key[149] = 6532890;
assign key2[149] = 9210;
assign key[150] = 6551300;
assign key2[150] = 9199;
assign key[151] = 6569688;
assign key2[151] = 9188;
assign key[152] = 6588053;
assign key2[152] = 9176;
assign key[153] = 6606395;
assign key2[153] = 9165;
assign key[154] = 6624716;
assign key2[154] = 9154;
assign key[155] = 6643013;
assign key2[155] = 9143;
assign key[156] = 6661289;
assign key2[156] = 9132;
assign key[157] = 6679542;
assign key2[157] = 9121;
assign key[158] = 6697774;
assign key2[158] = 9110;
assign key[159] = 6715983;
assign key2[159] = 9099;
assign key[160] = 6734170;
assign key2[160] = 9088;
assign key[161] = 6752336;
assign key2[161] = 9077;
assign key[162] = 6770479;
assign key2[162] = 9066;
assign key[163] = 6788601;
assign key2[163] = 9055;
assign key[164] = 6806702;
assign key2[164] = 9044;
assign key[165] = 6824781;
assign key2[165] = 9034;
assign key[166] = 6842838;
assign key2[166] = 9023;
assign key[167] = 6860874;
assign key2[167] = 9012;
assign key[168] = 6878889;
assign key2[168] = 9002;
assign key[169] = 6896883;
assign key2[169] = 8991;
assign key[170] = 6914855;
assign key2[170] = 8980;
assign key[171] = 6932806;
assign key2[171] = 8970;
assign key[172] = 6950736;
assign key2[172] = 8959;
assign key[173] = 6968646;
assign key2[173] = 8949;
assign key[174] = 6986534;
assign key2[174] = 8939;
assign key[175] = 7004402;
assign key2[175] = 8928;
assign key[176] = 7022249;
assign key2[176] = 8918;
assign key[177] = 7040075;
assign key2[177] = 8908;
assign key[178] = 7057881;
assign key2[178] = 8897;
assign key[179] = 7075666;
assign key2[179] = 8887;
assign key[180] = 7093431;
assign key2[180] = 8877;
assign key[181] = 7111176;
assign key2[181] = 8867;
assign key[182] = 7128900;
assign key2[182] = 8857;
assign key[183] = 7146604;
assign key2[183] = 8846;
assign key[184] = 7164287;
assign key2[184] = 8836;
assign key[185] = 7181951;
assign key2[185] = 8826;
assign key[186] = 7199595;
assign key2[186] = 8816;
assign key[187] = 7217219;
assign key2[187] = 8806;
assign key[188] = 7234823;
assign key2[188] = 8796;
assign key[189] = 7252407;
assign key2[189] = 8787;
assign key[190] = 7269971;
assign key2[190] = 8777;
assign key[191] = 7287516;
assign key2[191] = 8767;
assign key[192] = 7305041;
assign key2[192] = 8757;
assign key[193] = 7322546;
assign key2[193] = 8747;
assign key[194] = 7340032;
assign key2[194] = 8738;
assign key[195] = 7357499;
assign key2[195] = 8728;
assign key[196] = 7374946;
assign key2[196] = 8718;
assign key[197] = 7392374;
assign key2[197] = 8709;
assign key[198] = 7409782;
assign key2[198] = 8699;
assign key[199] = 7427172;
assign key2[199] = 8689;
assign key[200] = 7444542;
assign key2[200] = 8680;
assign key[201] = 7461894;
assign key2[201] = 8670;
assign key[202] = 7479226;
assign key2[202] = 8661;
assign key[203] = 7496540;
assign key2[203] = 8652;
assign key[204] = 7513834;
assign key2[204] = 8642;
assign key[205] = 7531110;
assign key2[205] = 8633;
assign key[206] = 7548367;
assign key2[206] = 8623;
assign key[207] = 7565606;
assign key2[207] = 8614;
assign key[208] = 7582826;
assign key2[208] = 8605;
assign key[209] = 7600027;
assign key2[209] = 8596;
assign key[210] = 7617210;
assign key2[210] = 8586;
assign key[211] = 7634374;
assign key2[211] = 8577;
assign key[212] = 7651520;
assign key2[212] = 8568;
assign key[213] = 7668648;
assign key2[213] = 8559;
assign key[214] = 7685758;
assign key2[214] = 8550;
assign key[215] = 7702849;
assign key2[215] = 8541;
assign key[216] = 7719922;
assign key2[216] = 8532;
assign key[217] = 7736977;
assign key2[217] = 8523;
assign key[218] = 7754014;
assign key2[218] = 8514;
assign key[219] = 7771033;
assign key2[219] = 8505;
assign key[220] = 7788035;
assign key2[220] = 8496;
assign key[221] = 7805018;
assign key2[221] = 8487;
assign key[222] = 7821984;
assign key2[222] = 8478;
assign key[223] = 7838931;
assign key2[223] = 8469;
assign key[224] = 7855862;
assign key2[224] = 8460;
assign key[225] = 7872774;
assign key2[225] = 8451;
assign key[226] = 7889669;
assign key2[226] = 8443;
assign key[227] = 7906546;
assign key2[227] = 8434;
assign key[228] = 7923406;
assign key2[228] = 8425;
assign key[229] = 7940249;
assign key2[229] = 8416;
assign key[230] = 7957074;
assign key2[230] = 8408;
assign key[231] = 7973882;
assign key2[231] = 8399;
assign key[232] = 7990673;
assign key2[232] = 8391;
assign key[233] = 8007446;
assign key2[233] = 8382;
assign key[234] = 8024203;
assign key2[234] = 8373;
assign key[235] = 8040942;
assign key2[235] = 8365;
assign key[236] = 8057664;
assign key2[236] = 8356;
assign key[237] = 8074369;
assign key2[237] = 8348;
assign key[238] = 8091057;
assign key2[238] = 8339;
assign key[239] = 8107729;
assign key2[239] = 8331;
assign key[240] = 8124383;
assign key2[240] = 8323;
assign key[241] = 8141021;
assign key2[241] = 8314;
assign key[242] = 8157642;
assign key2[242] = 8306;
assign key[243] = 8174247;
assign key2[243] = 8298;
assign key[244] = 8190834;
assign key2[244] = 8289;
assign key[245] = 8207405;
assign key2[245] = 8281;
assign key[246] = 8223960;
assign key2[246] = 8273;
assign key[247] = 8240498;
assign key2[247] = 8264;
assign key[248] = 8257020;
assign key2[248] = 8256;
assign key[249] = 8273525;
assign key2[249] = 8248;
assign key[250] = 8290014;
assign key2[250] = 8240;
assign key[251] = 8306487;
assign key2[251] = 8232;
assign key[252] = 8322943;
assign key2[252] = 8224;
assign key[253] = 8339384;
assign key2[253] = 8216;
assign key[254] = 8355808;
assign key2[254] = 8208;
assign key[255] = 8372216;
assign key2[255] = 8200;
assign key[256] = 0;
assign key2[256] = 8192;
assign key[257] = 16368;
assign key2[257] = 8176;
assign key[258] = 32704;
assign key2[258] = 8160;
assign key[259] = 49009;
assign key2[259] = 8144;
assign key[260] = 65282;
assign key2[260] = 8128;
assign key[261] = 81524;
assign key2[261] = 8113;
assign key[262] = 97735;
assign key2[262] = 8097;
assign key[263] = 113915;
assign key2[263] = 8082;
assign key[264] = 130064;
assign key2[264] = 8066;
assign key[265] = 146182;
assign key2[265] = 8051;
assign key[266] = 162271;
assign key2[266] = 8036;
assign key[267] = 178329;
assign key2[267] = 8021;
assign key[268] = 194356;
assign key2[268] = 8006;
assign key[269] = 210355;
assign key2[269] = 7991;
assign key[270] = 226323;
assign key2[270] = 7976;
assign key[271] = 242262;
assign key2[271] = 7962;
assign key[272] = 258171;
assign key2[272] = 7947;
assign key[273] = 274051;
assign key2[273] = 7932;
assign key[274] = 289903;
assign key2[274] = 7918;
assign key[275] = 305725;
assign key2[275] = 7903;
assign key[276] = 321518;
assign key2[276] = 7889;
assign key[277] = 337283;
assign key2[277] = 7875;
assign key[278] = 353020;
assign key2[278] = 7861;
assign key[279] = 368728;
assign key2[279] = 7847;
assign key[280] = 384408;
assign key2[280] = 7833;
assign key[281] = 400060;
assign key2[281] = 7819;
assign key[282] = 415685;
assign key2[282] = 7805;
assign key[283] = 431281;
assign key2[283] = 7791;
assign key[284] = 446850;
assign key2[284] = 7777;
assign key[285] = 462392;
assign key2[285] = 7764;
assign key[286] = 477907;
assign key2[286] = 7750;
assign key[287] = 493394;
assign key2[287] = 7736;
assign key[288] = 508854;
assign key2[288] = 7723;
assign key[289] = 524288;
assign key2[289] = 7710;
assign key[290] = 539695;
assign key2[290] = 7696;
assign key[291] = 555075;
assign key2[291] = 7683;
assign key[292] = 570429;
assign key2[292] = 7670;
assign key[293] = 585757;
assign key2[293] = 7657;
assign key[294] = 601059;
assign key2[294] = 7644;
assign key[295] = 616334;
assign key2[295] = 7631;
assign key[296] = 631584;
assign key2[296] = 7618;
assign key[297] = 646808;
assign key2[297] = 7605;
assign key[298] = 662006;
assign key2[298] = 7592;
assign key[299] = 677179;
assign key2[299] = 7580;
assign key[300] = 692327;
assign key2[300] = 7567;
assign key[301] = 707449;
assign key2[301] = 7554;
assign key[302] = 722546;
assign key2[302] = 7542;
assign key[303] = 737618;
assign key2[303] = 7529;
assign key[304] = 752666;
assign key2[304] = 7517;
assign key[305] = 767688;
assign key2[305] = 7505;
assign key[306] = 782686;
assign key2[306] = 7492;
assign key[307] = 797660;
assign key2[307] = 7480;
assign key[308] = 812609;
assign key2[308] = 7468;
assign key[309] = 827534;
assign key2[309] = 7456;
assign key[310] = 842435;
assign key2[310] = 7444;
assign key[311] = 857312;
assign key2[311] = 7432;
assign key[312] = 872164;
assign key2[312] = 7420;
assign key[313] = 886994;
assign key2[313] = 7408;
assign key[314] = 901799;
assign key2[314] = 7396;
assign key[315] = 916581;
assign key2[315] = 7385;
assign key[316] = 931339;
assign key2[316] = 7373;
assign key[317] = 946074;
assign key2[317] = 7361;
assign key[318] = 960786;
assign key2[318] = 7350;
assign key[319] = 975475;
assign key2[319] = 7338;
assign key[320] = 990141;
assign key2[320] = 7327;
assign key[321] = 1004784;
assign key2[321] = 7315;
assign key[322] = 1019404;
assign key2[322] = 7304;
assign key[323] = 1034001;
assign key2[323] = 7293;
assign key[324] = 1048576;
assign key2[324] = 7281;
assign key[325] = 1063128;
assign key2[325] = 7270;
assign key[326] = 1077658;
assign key2[326] = 7259;
assign key[327] = 1092166;
assign key2[327] = 7248;
assign key[328] = 1106652;
assign key2[328] = 7237;
assign key[329] = 1121115;
assign key2[329] = 7226;
assign key[330] = 1135556;
assign key2[330] = 7215;
assign key[331] = 1149976;
assign key2[331] = 7204;
assign key[332] = 1164374;
assign key2[332] = 7193;
assign key[333] = 1178750;
assign key2[333] = 7182;
assign key[334] = 1193105;
assign key2[334] = 7171;
assign key[335] = 1207438;
assign key2[335] = 7161;
assign key[336] = 1221750;
assign key2[336] = 7150;
assign key[337] = 1236040;
assign key2[337] = 7139;
assign key[338] = 1250310;
assign key2[338] = 7129;
assign key[339] = 1264558;
assign key2[339] = 7118;
assign key[340] = 1278785;
assign key2[340] = 7108;
assign key[341] = 1292991;
assign key2[341] = 7097;
assign key[342] = 1307177;
assign key2[342] = 7087;
assign key[343] = 1321342;
assign key2[343] = 7077;
assign key[344] = 1335486;
assign key2[344] = 7066;
assign key[345] = 1349609;
assign key2[345] = 7056;
assign key[346] = 1363713;
assign key2[346] = 7046;
assign key[347] = 1377795;
assign key2[347] = 7036;
assign key[348] = 1391858;
assign key2[348] = 7026;
assign key[349] = 1405900;
assign key2[349] = 7016;
assign key[350] = 1419922;
assign key2[350] = 7006;
assign key[351] = 1433925;
assign key2[351] = 6996;
assign key[352] = 1447907;
assign key2[352] = 6986;
assign key[353] = 1461869;
assign key2[353] = 6976;
assign key[354] = 1475812;
assign key2[354] = 6966;
assign key[355] = 1489735;
assign key2[355] = 6956;
assign key[356] = 1503638;
assign key2[356] = 6946;
assign key[357] = 1517522;
assign key2[357] = 6937;
assign key[358] = 1531386;
assign key2[358] = 6927;
assign key[359] = 1545232;
assign key2[359] = 6917;
assign key[360] = 1559057;
assign key2[360] = 6908;
assign key[361] = 1572864;
assign key2[361] = 6898;
assign key[362] = 1586652;
assign key2[362] = 6888;
assign key[363] = 1600420;
assign key2[363] = 6879;
assign key[364] = 1614170;
assign key2[364] = 6870;
assign key[365] = 1627900;
assign key2[365] = 6860;
assign key[366] = 1641612;
assign key2[366] = 6851;
assign key[367] = 1655305;
assign key2[367] = 6841;
assign key[368] = 1668980;
assign key2[368] = 6832;
assign key[369] = 1682636;
assign key2[369] = 6823;
assign key[370] = 1696273;
assign key2[370] = 6814;
assign key[371] = 1709892;
assign key2[371] = 6804;
assign key[372] = 1723493;
assign key2[372] = 6795;
assign key[373] = 1737075;
assign key2[373] = 6786;
assign key[374] = 1750639;
assign key2[374] = 6777;
assign key[375] = 1764185;
assign key2[375] = 6768;
assign key[376] = 1777714;
assign key2[376] = 6759;
assign key[377] = 1791224;
assign key2[377] = 6750;
assign key[378] = 1804716;
assign key2[378] = 6741;
assign key[379] = 1818190;
assign key2[379] = 6732;
assign key[380] = 1831647;
assign key2[380] = 6723;
assign key[381] = 1845085;
assign key2[381] = 6715;
assign key[382] = 1858507;
assign key2[382] = 6706;
assign key[383] = 1871910;
assign key2[383] = 6697;
assign key[384] = 1885297;
assign key2[384] = 6688;
assign key[385] = 1898665;
assign key2[385] = 6680;
assign key[386] = 1912017;
assign key2[386] = 6671;
assign key[387] = 1925351;
assign key2[387] = 6662;
assign key[388] = 1938668;
assign key2[388] = 6654;
assign key[389] = 1951968;
assign key2[389] = 6645;
assign key[390] = 1965250;
assign key2[390] = 6637;
assign key[391] = 1978516;
assign key2[391] = 6628;
assign key[392] = 1991765;
assign key2[392] = 6620;
assign key[393] = 2004997;
assign key2[393] = 6611;
assign key[394] = 2018212;
assign key2[394] = 6603;
assign key[395] = 2031410;
assign key2[395] = 6594;
assign key[396] = 2044591;
assign key2[396] = 6586;
assign key[397] = 2057756;
assign key2[397] = 6578;
assign key[398] = 2070905;
assign key2[398] = 6570;
assign key[399] = 2084037;
assign key2[399] = 6561;
assign key[400] = 2097152;
assign key2[400] = 6553;
assign key[401] = 2110251;
assign key2[401] = 6545;
assign key[402] = 2123334;
assign key2[402] = 6537;
assign key[403] = 2136400;
assign key2[403] = 6529;
assign key[404] = 2149450;
assign key2[404] = 6521;
assign key[405] = 2162484;
assign key2[405] = 6513;
assign key[406] = 2175502;
assign key2[406] = 6504;
assign key[407] = 2188504;
assign key2[407] = 6496;
assign key[408] = 2201490;
assign key2[408] = 6489;
assign key[409] = 2214461;
assign key2[409] = 6481;
assign key[410] = 2227415;
assign key2[410] = 6473;
assign key[411] = 2240353;
assign key2[411] = 6465;
assign key[412] = 2253276;
assign key2[412] = 6457;
assign key[413] = 2266183;
assign key2[413] = 6449;
assign key[414] = 2279075;
assign key2[414] = 6441;
assign key[415] = 2291951;
assign key2[415] = 6434;
assign key[416] = 2304811;
assign key2[416] = 6426;
assign key[417] = 2317656;
assign key2[417] = 6418;
assign key[418] = 2330485;
assign key2[418] = 6410;
assign key[419] = 2343300;
assign key2[419] = 6403;
assign key[420] = 2356099;
assign key2[420] = 6395;
assign key[421] = 2368882;
assign key2[421] = 6388;
assign key[422] = 2381651;
assign key2[422] = 6380;
assign key[423] = 2394404;
assign key2[423] = 6372;
assign key[424] = 2407143;
assign key2[424] = 6365;
assign key[425] = 2419866;
assign key2[425] = 6357;
assign key[426] = 2432574;
assign key2[426] = 6350;
assign key[427] = 2445268;
assign key2[427] = 6343;
assign key[428] = 2457946;
assign key2[428] = 6335;
assign key[429] = 2470610;
assign key2[429] = 6328;
assign key[430] = 2483259;
assign key2[430] = 6320;
assign key[431] = 2495894;
assign key2[431] = 6313;
assign key[432] = 2508513;
assign key2[432] = 6306;
assign key[433] = 2521119;
assign key2[433] = 6298;
assign key[434] = 2533709;
assign key2[434] = 6291;
assign key[435] = 2546285;
assign key2[435] = 6284;
assign key[436] = 2558847;
assign key2[436] = 6277;
assign key[437] = 2571394;
assign key2[437] = 6270;
assign key[438] = 2583927;
assign key2[438] = 6262;
assign key[439] = 2596446;
assign key2[439] = 6255;
assign key[440] = 2608950;
assign key2[440] = 6248;
assign key[441] = 2621440;
assign key2[441] = 6241;
assign key[442] = 2633916;
assign key2[442] = 6234;
assign key[443] = 2646378;
assign key2[443] = 6227;
assign key[444] = 2658826;
assign key2[444] = 6220;
assign key[445] = 2671259;
assign key2[445] = 6213;
assign key[446] = 2683679;
assign key2[446] = 6206;
assign key[447] = 2696085;
assign key2[447] = 6199;
assign key[448] = 2708477;
assign key2[448] = 6192;
assign key[449] = 2720856;
assign key2[449] = 6185;
assign key[450] = 2733220;
assign key2[450] = 6178;
assign key[451] = 2745571;
assign key2[451] = 6171;
assign key[452] = 2757908;
assign key2[452] = 6165;
assign key[453] = 2770231;
assign key2[453] = 6158;
assign key[454] = 2782541;
assign key2[454] = 6151;
assign key[455] = 2794837;
assign key2[455] = 6144;
assign key[456] = 2807120;
assign key2[456] = 6138;
assign key[457] = 2819389;
assign key2[457] = 6131;
assign key[458] = 2831645;
assign key2[458] = 6124;
assign key[459] = 2843888;
assign key2[459] = 6117;
assign key[460] = 2856117;
assign key2[460] = 6111;
assign key[461] = 2868333;
assign key2[461] = 6104;
assign key[462] = 2880535;
assign key2[462] = 6098;
assign key[463] = 2892725;
assign key2[463] = 6091;
assign key[464] = 2904901;
assign key2[464] = 6084;
assign key[465] = 2917064;
assign key2[465] = 6078;
assign key[466] = 2929214;
assign key2[466] = 6071;
assign key[467] = 2941352;
assign key2[467] = 6065;
assign key[468] = 2953476;
assign key2[468] = 6058;
assign key[469] = 2965587;
assign key2[469] = 6052;
assign key[470] = 2977685;
assign key2[470] = 6045;
assign key[471] = 2989770;
assign key2[471] = 6039;
assign key[472] = 3001843;
assign key2[472] = 6033;
assign key[473] = 3013903;
assign key2[473] = 6026;
assign key[474] = 3025950;
assign key2[474] = 6020;
assign key[475] = 3037984;
assign key2[475] = 6013;
assign key[476] = 3050006;
assign key2[476] = 6007;
assign key[477] = 3062015;
assign key2[477] = 6001;
assign key[478] = 3074011;
assign key2[478] = 5995;
assign key[479] = 3085995;
assign key2[479] = 5988;
assign key[480] = 3097967;
assign key2[480] = 5982;
assign key[481] = 3109926;
assign key2[481] = 5976;
assign key[482] = 3121872;
assign key2[482] = 5970;
assign key[483] = 3133806;
assign key2[483] = 5963;
assign key[484] = 3145728;
assign key2[484] = 5957;
assign key[485] = 3157637;
assign key2[485] = 5951;
assign key[486] = 3169535;
assign key2[486] = 5945;
assign key[487] = 3181420;
assign key2[487] = 5939;
assign key[488] = 3193292;
assign key2[488] = 5933;
assign key[489] = 3205153;
assign key2[489] = 5927;
assign key[490] = 3217002;
assign key2[490] = 5921;
assign key[491] = 3228838;
assign key2[491] = 5915;
assign key[492] = 3240662;
assign key2[492] = 5909;
assign key[493] = 3252475;
assign key2[493] = 5903;
assign key[494] = 3264275;
assign key2[494] = 5897;
assign key[495] = 3276064;
assign key2[495] = 5891;
assign key[496] = 3287840;
assign key2[496] = 5885;
assign key[497] = 3299605;
assign key2[497] = 5879;
assign key[498] = 3311358;
assign key2[498] = 5873;
assign key[499] = 3323099;
assign key2[499] = 5867;
assign key[500] = 3334828;
assign key2[500] = 5861;
assign key[501] = 3346546;
assign key2[501] = 5855;
assign key[502] = 3358252;
assign key2[502] = 5850;
assign key[503] = 3369946;
assign key2[503] = 5844;
assign key[504] = 3381628;
assign key2[504] = 5838;
assign key[505] = 3393299;
assign key2[505] = 5832;
assign key[506] = 3404959;
assign key2[506] = 5826;
assign key[507] = 3416607;
assign key2[507] = 5821;
assign key[508] = 3428243;
assign key2[508] = 5815;
assign key[509] = 3439868;
assign key2[509] = 5809;
assign key[510] = 3451482;
assign key2[510] = 5803;
assign key[511] = 3463084;
assign key2[511] = 5798;

wire [8:0] se;
assign se = adata[23] ? {1'b0,((adata[30:23] >> 1) + 8'd64)} : {1'b0,((adata[30:23] >> 1) + 8'd63)};

wire [8:0] index;
assign index = adata[23:15];

/*
wire [14:0] b;
assign b = adata[14] ? ~adata[14:0]+1 : adata[14:0];

wire [13:0] k;
assign k = adata[14] ? key2[index+1] : key2[index];
*/

wire [22:0] a;
assign a = adata[14] ? key[index+1] : key[index];

wire check;
assign check = ~(|(~adata[22:14]));

/*
wire [28:0] bk;
assign bk = b * k;
*/

wire [14:0] kuso;
assign kuso = ~adata[14:0]+15'b1;

wire [28:0] bkxk;
assign bkxk = kuso * 5792;

wire [28:0] bkxg;
assign bkxg = kuso * 8192;

wire [28:0] bkn;
assign bkn = kuso * key2[index+1];

wire [28:0] bkp;
assign bkp = adata[14:0] * key2[index];


reg [22:0] a_reg;
reg check_reg;
reg [28:0] bkxk_reg;
reg [28:0] bkxg_reg;
reg [28:0] bkn_reg;
reg [28:0] bkp_reg;
reg notzero_reg;
reg [8:0] se_reg;
reg adata14_reg;
reg adata23_reg;
reg flag_reg;
reg [4:0] address_reg;

always_ff@(posedge clk) begin
a_reg <= check ? (adata[23] ? 3474675 : 8388607) : a;
check_reg <= check;
bkxk_reg <= bkxk;
bkxg_reg <= bkxg;
bkn_reg <= bkn;
bkp_reg <= bkp; 
notzero_reg <= |adata[30:23];
se_reg <= se;
adata14_reg <= adata[14];
adata23_reg <= adata[23];
flag_reg <= flag_in;
address_reg <= address_in;
end


/*
wire [22:0] a_reg;
wire [28:0] bk_reg;
wire notzero_reg;
wire [8:0] se_reg;
wire adata14_reg;
wire flag_reg;
wire [4:0] address_reg;

assign a_reg = check ? (adata[23] ? 3474675 : 8388607) : a;
assign bk_reg = check ? bkx : bk;
assign notzero_reg = |adata[30:23];
assign se_reg = se;
assign adata14_reg = adata[14];
assign flag_reg = flag_in;
assign address_reg = address_in;

*/

wire [28:0] bk;
assign bk = check_reg ? (adata23_reg ? bkxk_reg : bkxg_reg) : (adata14_reg ? bkn_reg : bkp_reg);

wire [14:0] bk2;
assign bk2 = bk[28:14];

wire [22:0] kari;
assign kari = adata14_reg ? a_reg - bk2 : a_reg + bk2;



always_ff@(posedge clk) begin
result <= notzero_reg ? {se_reg,kari} : 0;
flag_out <= flag_reg;
address_out <= address_reg;
end

endmodule

`default_nettype wire
