`default_nettype none

module fdiv(
input wire [31:0] adata,
input wire [31:0] bdata,
output reg [31:0] result,
input wire clk,
input wire flag_in,
input wire [4:0] address_in,
output reg flag_out,
output reg [4:0] address_out);

reg [24:0] s [2047:0];
reg [12:0] t [2047:0];

assign s[0] = 16777216;
assign t[0] = 8188;
assign s[1] = 16769028;
assign t[1] = 8180;
assign s[2] = 16760847;
assign t[2] = 8172;
assign s[3] = 16752675;
assign t[3] = 8164;
assign s[4] = 16744511;
assign t[4] = 8156;
assign s[5] = 16736355;
assign t[5] = 8148;
assign s[6] = 16728207;
assign t[6] = 8140;
assign s[7] = 16720067;
assign t[7] = 8132;
assign s[8] = 16711935;
assign t[8] = 8124;
assign s[9] = 16703810;
assign t[9] = 8116;
assign s[10] = 16695694;
assign t[10] = 8108;
assign s[11] = 16687585;
assign t[11] = 8100;
assign s[12] = 16679484;
assign t[12] = 8092;
assign s[13] = 16671391;
assign t[13] = 8085;
assign s[14] = 16663306;
assign t[14] = 8077;
assign s[15] = 16655229;
assign t[15] = 8069;
assign s[16] = 16647160;
assign t[16] = 8061;
assign s[17] = 16639098;
assign t[17] = 8053;
assign s[18] = 16631044;
assign t[18] = 8045;
assign s[19] = 16622998;
assign t[19] = 8038;
assign s[20] = 16614960;
assign t[20] = 8030;
assign s[21] = 16606930;
assign t[21] = 8022;
assign s[22] = 16598907;
assign t[22] = 8014;
assign s[23] = 16590892;
assign t[23] = 8007;
assign s[24] = 16582885;
assign t[24] = 7999;
assign s[25] = 16574885;
assign t[25] = 7991;
assign s[26] = 16566894;
assign t[26] = 7984;
assign s[27] = 16558910;
assign t[27] = 7976;
assign s[28] = 16550933;
assign t[28] = 7968;
assign s[29] = 16542965;
assign t[29] = 7961;
assign s[30] = 16535004;
assign t[30] = 7953;
assign s[31] = 16527050;
assign t[31] = 7945;
assign s[32] = 16519105;
assign t[32] = 7938;
assign s[33] = 16511166;
assign t[33] = 7930;
assign s[34] = 16503236;
assign t[34] = 7922;
assign s[35] = 16495313;
assign t[35] = 7915;
assign s[36] = 16487398;
assign t[36] = 7907;
assign s[37] = 16479490;
assign t[37] = 7900;
assign s[38] = 16471590;
assign t[38] = 7892;
assign s[39] = 16463698;
assign t[39] = 7884;
assign s[40] = 16455813;
assign t[40] = 7877;
assign s[41] = 16447936;
assign t[41] = 7869;
assign s[42] = 16440066;
assign t[42] = 7862;
assign s[43] = 16432203;
assign t[43] = 7854;
assign s[44] = 16424349;
assign t[44] = 7847;
assign s[45] = 16416501;
assign t[45] = 7839;
assign s[46] = 16408662;
assign t[46] = 7832;
assign s[47] = 16400829;
assign t[47] = 7824;
assign s[48] = 16393005;
assign t[48] = 7817;
assign s[49] = 16385187;
assign t[49] = 7809;
assign s[50] = 16377377;
assign t[50] = 7802;
assign s[51] = 16369575;
assign t[51] = 7795;
assign s[52] = 16361780;
assign t[52] = 7787;
assign s[53] = 16353992;
assign t[53] = 7780;
assign s[54] = 16346212;
assign t[54] = 7772;
assign s[55] = 16338439;
assign t[55] = 7765;
assign s[56] = 16330674;
assign t[56] = 7758;
assign s[57] = 16322916;
assign t[57] = 7750;
assign s[58] = 16315165;
assign t[58] = 7743;
assign s[59] = 16307422;
assign t[59] = 7735;
assign s[60] = 16299686;
assign t[60] = 7728;
assign s[61] = 16291957;
assign t[61] = 7721;
assign s[62] = 16284236;
assign t[62] = 7713;
assign s[63] = 16276522;
assign t[63] = 7706;
assign s[64] = 16268815;
assign t[64] = 7699;
assign s[65] = 16261116;
assign t[65] = 7692;
assign s[66] = 16253424;
assign t[66] = 7684;
assign s[67] = 16245739;
assign t[67] = 7677;
assign s[68] = 16238061;
assign t[68] = 7670;
assign s[69] = 16230391;
assign t[69] = 7663;
assign s[70] = 16222728;
assign t[70] = 7655;
assign s[71] = 16215072;
assign t[71] = 7648;
assign s[72] = 16207423;
assign t[72] = 7641;
assign s[73] = 16199782;
assign t[73] = 7634;
assign s[74] = 16192148;
assign t[74] = 7627;
assign s[75] = 16184521;
assign t[75] = 7619;
assign s[76] = 16176901;
assign t[76] = 7612;
assign s[77] = 16169288;
assign t[77] = 7605;
assign s[78] = 16161683;
assign t[78] = 7598;
assign s[79] = 16154084;
assign t[79] = 7591;
assign s[80] = 16146493;
assign t[80] = 7584;
assign s[81] = 16138909;
assign t[81] = 7576;
assign s[82] = 16131332;
assign t[82] = 7569;
assign s[83] = 16123762;
assign t[83] = 7562;
assign s[84] = 16116200;
assign t[84] = 7555;
assign s[85] = 16108644;
assign t[85] = 7548;
assign s[86] = 16101095;
assign t[86] = 7541;
assign s[87] = 16093554;
assign t[87] = 7534;
assign s[88] = 16086019;
assign t[88] = 7527;
assign s[89] = 16078492;
assign t[89] = 7520;
assign s[90] = 16070972;
assign t[90] = 7513;
assign s[91] = 16063458;
assign t[91] = 7506;
assign s[92] = 16055952;
assign t[92] = 7499;
assign s[93] = 16048453;
assign t[93] = 7492;
assign s[94] = 16040961;
assign t[94] = 7485;
assign s[95] = 16033475;
assign t[95] = 7478;
assign s[96] = 16025997;
assign t[96] = 7471;
assign s[97] = 16018526;
assign t[97] = 7464;
assign s[98] = 16011061;
assign t[98] = 7457;
assign s[99] = 16003604;
assign t[99] = 7450;
assign s[100] = 15996153;
assign t[100] = 7443;
assign s[101] = 15988710;
assign t[101] = 7436;
assign s[102] = 15981273;
assign t[102] = 7429;
assign s[103] = 15973844;
assign t[103] = 7422;
assign s[104] = 15966421;
assign t[104] = 7415;
assign s[105] = 15959005;
assign t[105] = 7409;
assign s[106] = 15951596;
assign t[106] = 7402;
assign s[107] = 15944194;
assign t[107] = 7395;
assign s[108] = 15936799;
assign t[108] = 7388;
assign s[109] = 15929410;
assign t[109] = 7381;
assign s[110] = 15922029;
assign t[110] = 7374;
assign s[111] = 15914654;
assign t[111] = 7367;
assign s[112] = 15907286;
assign t[112] = 7361;
assign s[113] = 15899925;
assign t[113] = 7354;
assign s[114] = 15892571;
assign t[114] = 7347;
assign s[115] = 15885223;
assign t[115] = 7340;
assign s[116] = 15877882;
assign t[116] = 7333;
assign s[117] = 15870549;
assign t[117] = 7327;
assign s[118] = 15863221;
assign t[118] = 7320;
assign s[119] = 15855901;
assign t[119] = 7313;
assign s[120] = 15848587;
assign t[120] = 7306;
assign s[121] = 15841281;
assign t[121] = 7300;
assign s[122] = 15833980;
assign t[122] = 7293;
assign s[123] = 15826687;
assign t[123] = 7286;
assign s[124] = 15819400;
assign t[124] = 7279;
assign s[125] = 15812120;
assign t[125] = 7273;
assign s[126] = 15804847;
assign t[126] = 7266;
assign s[127] = 15797581;
assign t[127] = 7259;
assign s[128] = 15790321;
assign t[128] = 7253;
assign s[129] = 15783067;
assign t[129] = 7246;
assign s[130] = 15775821;
assign t[130] = 7239;
assign s[131] = 15768581;
assign t[131] = 7233;
assign s[132] = 15761348;
assign t[132] = 7226;
assign s[133] = 15754121;
assign t[133] = 7220;
assign s[134] = 15746901;
assign t[134] = 7213;
assign s[135] = 15739687;
assign t[135] = 7206;
assign s[136] = 15732481;
assign t[136] = 7200;
assign s[137] = 15725280;
assign t[137] = 7193;
assign s[138] = 15718087;
assign t[138] = 7187;
assign s[139] = 15710900;
assign t[139] = 7180;
assign s[140] = 15703719;
assign t[140] = 7173;
assign s[141] = 15696545;
assign t[141] = 7167;
assign s[142] = 15689378;
assign t[142] = 7160;
assign s[143] = 15682217;
assign t[143] = 7154;
assign s[144] = 15675063;
assign t[144] = 7147;
assign s[145] = 15667915;
assign t[145] = 7141;
assign s[146] = 15660774;
assign t[146] = 7134;
assign s[147] = 15653639;
assign t[147] = 7128;
assign s[148] = 15646511;
assign t[148] = 7121;
assign s[149] = 15639389;
assign t[149] = 7115;
assign s[150] = 15632274;
assign t[150] = 7108;
assign s[151] = 15625165;
assign t[151] = 7102;
assign s[152] = 15618063;
assign t[152] = 7095;
assign s[153] = 15610967;
assign t[153] = 7089;
assign s[154] = 15603877;
assign t[154] = 7083;
assign s[155] = 15596794;
assign t[155] = 7076;
assign s[156] = 15589718;
assign t[156] = 7070;
assign s[157] = 15582647;
assign t[157] = 7063;
assign s[158] = 15575584;
assign t[158] = 7057;
assign s[159] = 15568526;
assign t[159] = 7050;
assign s[160] = 15561475;
assign t[160] = 7044;
assign s[161] = 15554431;
assign t[161] = 7038;
assign s[162] = 15547393;
assign t[162] = 7031;
assign s[163] = 15540361;
assign t[163] = 7025;
assign s[164] = 15533335;
assign t[164] = 7019;
assign s[165] = 15526316;
assign t[165] = 7012;
assign s[166] = 15519303;
assign t[166] = 7006;
assign s[167] = 15512297;
assign t[167] = 7000;
assign s[168] = 15505297;
assign t[168] = 6993;
assign s[169] = 15498303;
assign t[169] = 6987;
assign s[170] = 15491315;
assign t[170] = 6981;
assign s[171] = 15484334;
assign t[171] = 6974;
assign s[172] = 15477359;
assign t[172] = 6968;
assign s[173] = 15470391;
assign t[173] = 6962;
assign s[174] = 15463428;
assign t[174] = 6956;
assign s[175] = 15456472;
assign t[175] = 6949;
assign s[176] = 15449522;
assign t[176] = 6943;
assign s[177] = 15442579;
assign t[177] = 6937;
assign s[178] = 15435641;
assign t[178] = 6931;
assign s[179] = 15428710;
assign t[179] = 6924;
assign s[180] = 15421785;
assign t[180] = 6918;
assign s[181] = 15414867;
assign t[181] = 6912;
assign s[182] = 15407954;
assign t[182] = 6906;
assign s[183] = 15401048;
assign t[183] = 6900;
assign s[184] = 15394148;
assign t[184] = 6893;
assign s[185] = 15387254;
assign t[185] = 6887;
assign s[186] = 15380366;
assign t[186] = 6881;
assign s[187] = 15373484;
assign t[187] = 6875;
assign s[188] = 15366609;
assign t[188] = 6869;
assign s[189] = 15359740;
assign t[189] = 6863;
assign s[190] = 15352877;
assign t[190] = 6857;
assign s[191] = 15346020;
assign t[191] = 6850;
assign s[192] = 15339169;
assign t[192] = 6844;
assign s[193] = 15332324;
assign t[193] = 6838;
assign s[194] = 15325485;
assign t[194] = 6832;
assign s[195] = 15318653;
assign t[195] = 6826;
assign s[196] = 15311826;
assign t[196] = 6820;
assign s[197] = 15305006;
assign t[197] = 6814;
assign s[198] = 15298191;
assign t[198] = 6808;
assign s[199] = 15291383;
assign t[199] = 6802;
assign s[200] = 15284581;
assign t[200] = 6796;
assign s[201] = 15277785;
assign t[201] = 6790;
assign s[202] = 15270995;
assign t[202] = 6784;
assign s[203] = 15264210;
assign t[203] = 6778;
assign s[204] = 15257432;
assign t[204] = 6772;
assign s[205] = 15250660;
assign t[205] = 6766;
assign s[206] = 15243894;
assign t[206] = 6760;
assign s[207] = 15237134;
assign t[207] = 6754;
assign s[208] = 15230380;
assign t[208] = 6748;
assign s[209] = 15223632;
assign t[209] = 6742;
assign s[210] = 15216890;
assign t[210] = 6736;
assign s[211] = 15210154;
assign t[211] = 6730;
assign s[212] = 15203424;
assign t[212] = 6724;
assign s[213] = 15196700;
assign t[213] = 6718;
assign s[214] = 15189981;
assign t[214] = 6712;
assign s[215] = 15183269;
assign t[215] = 6706;
assign s[216] = 15176563;
assign t[216] = 6700;
assign s[217] = 15169862;
assign t[217] = 6694;
assign s[218] = 15163168;
assign t[218] = 6688;
assign s[219] = 15156479;
assign t[219] = 6682;
assign s[220] = 15149796;
assign t[220] = 6676;
assign s[221] = 15143119;
assign t[221] = 6670;
assign s[222] = 15136448;
assign t[222] = 6665;
assign s[223] = 15129783;
assign t[223] = 6659;
assign s[224] = 15123124;
assign t[224] = 6653;
assign s[225] = 15116471;
assign t[225] = 6647;
assign s[226] = 15109823;
assign t[226] = 6641;
assign s[227] = 15103181;
assign t[227] = 6635;
assign s[228] = 15096546;
assign t[228] = 6630;
assign s[229] = 15089916;
assign t[229] = 6624;
assign s[230] = 15083291;
assign t[230] = 6618;
assign s[231] = 15076673;
assign t[231] = 6612;
assign s[232] = 15070060;
assign t[232] = 6606;
assign s[233] = 15063454;
assign t[233] = 6600;
assign s[234] = 15056853;
assign t[234] = 6595;
assign s[235] = 15050257;
assign t[235] = 6589;
assign s[236] = 15043668;
assign t[236] = 6583;
assign s[237] = 15037084;
assign t[237] = 6577;
assign s[238] = 15030507;
assign t[238] = 6572;
assign s[239] = 15023934;
assign t[239] = 6566;
assign s[240] = 15017368;
assign t[240] = 6560;
assign s[241] = 15010807;
assign t[241] = 6554;
assign s[242] = 15004252;
assign t[242] = 6549;
assign s[243] = 14997703;
assign t[243] = 6543;
assign s[244] = 14991160;
assign t[244] = 6537;
assign s[245] = 14984622;
assign t[245] = 6532;
assign s[246] = 14978090;
assign t[246] = 6526;
assign s[247] = 14971563;
assign t[247] = 6520;
assign s[248] = 14965043;
assign t[248] = 6515;
assign s[249] = 14958528;
assign t[249] = 6509;
assign s[250] = 14952018;
assign t[250] = 6503;
assign s[251] = 14945515;
assign t[251] = 6498;
assign s[252] = 14939016;
assign t[252] = 6492;
assign s[253] = 14932524;
assign t[253] = 6486;
assign s[254] = 14926037;
assign t[254] = 6481;
assign s[255] = 14919556;
assign t[255] = 6475;
assign s[256] = 14913081;
assign t[256] = 6469;
assign s[257] = 14906611;
assign t[257] = 6464;
assign s[258] = 14900147;
assign t[258] = 6458;
assign s[259] = 14893688;
assign t[259] = 6453;
assign s[260] = 14887235;
assign t[260] = 6447;
assign s[261] = 14880787;
assign t[261] = 6441;
assign s[262] = 14874345;
assign t[262] = 6436;
assign s[263] = 14867909;
assign t[263] = 6430;
assign s[264] = 14861478;
assign t[264] = 6425;
assign s[265] = 14855053;
assign t[265] = 6419;
assign s[266] = 14848634;
assign t[266] = 6414;
assign s[267] = 14842219;
assign t[267] = 6408;
assign s[268] = 14835811;
assign t[268] = 6403;
assign s[269] = 14829408;
assign t[269] = 6397;
assign s[270] = 14823010;
assign t[270] = 6391;
assign s[271] = 14816618;
assign t[271] = 6386;
assign s[272] = 14810232;
assign t[272] = 6380;
assign s[273] = 14803851;
assign t[273] = 6375;
assign s[274] = 14797475;
assign t[274] = 6369;
assign s[275] = 14791105;
assign t[275] = 6364;
assign s[276] = 14784741;
assign t[276] = 6359;
assign s[277] = 14778382;
assign t[277] = 6353;
assign s[278] = 14772028;
assign t[278] = 6348;
assign s[279] = 14765680;
assign t[279] = 6342;
assign s[280] = 14759338;
assign t[280] = 6337;
assign s[281] = 14753000;
assign t[281] = 6331;
assign s[282] = 14746669;
assign t[282] = 6326;
assign s[283] = 14740342;
assign t[283] = 6320;
assign s[284] = 14734021;
assign t[284] = 6315;
assign s[285] = 14727706;
assign t[285] = 6310;
assign s[286] = 14721396;
assign t[286] = 6304;
assign s[287] = 14715091;
assign t[287] = 6299;
assign s[288] = 14708792;
assign t[288] = 6293;
assign s[289] = 14702498;
assign t[289] = 6288;
assign s[290] = 14696210;
assign t[290] = 6283;
assign s[291] = 14689926;
assign t[291] = 6277;
assign s[292] = 14683649;
assign t[292] = 6272;
assign s[293] = 14677376;
assign t[293] = 6267;
assign s[294] = 14671109;
assign t[294] = 6261;
assign s[295] = 14664848;
assign t[295] = 6256;
assign s[296] = 14658591;
assign t[296] = 6250;
assign s[297] = 14652340;
assign t[297] = 6245;
assign s[298] = 14646095;
assign t[298] = 6240;
assign s[299] = 14639854;
assign t[299] = 6235;
assign s[300] = 14633619;
assign t[300] = 6229;
assign s[301] = 14627390;
assign t[301] = 6224;
assign s[302] = 14621165;
assign t[302] = 6219;
assign s[303] = 14614946;
assign t[303] = 6213;
assign s[304] = 14608732;
assign t[304] = 6208;
assign s[305] = 14602524;
assign t[305] = 6203;
assign s[306] = 14596320;
assign t[306] = 6198;
assign s[307] = 14590122;
assign t[307] = 6192;
assign s[308] = 14583930;
assign t[308] = 6187;
assign s[309] = 14577742;
assign t[309] = 6182;
assign s[310] = 14571560;
assign t[310] = 6177;
assign s[311] = 14565383;
assign t[311] = 6171;
assign s[312] = 14559211;
assign t[312] = 6166;
assign s[313] = 14553044;
assign t[313] = 6161;
assign s[314] = 14546883;
assign t[314] = 6156;
assign s[315] = 14540727;
assign t[315] = 6150;
assign s[316] = 14534576;
assign t[316] = 6145;
assign s[317] = 14528430;
assign t[317] = 6140;
assign s[318] = 14522290;
assign t[318] = 6135;
assign s[319] = 14516155;
assign t[319] = 6130;
assign s[320] = 14510025;
assign t[320] = 6124;
assign s[321] = 14503900;
assign t[321] = 6119;
assign s[322] = 14497780;
assign t[322] = 6114;
assign s[323] = 14491665;
assign t[323] = 6109;
assign s[324] = 14485556;
assign t[324] = 6104;
assign s[325] = 14479451;
assign t[325] = 6099;
assign s[326] = 14473352;
assign t[326] = 6094;
assign s[327] = 14467258;
assign t[327] = 6088;
assign s[328] = 14461169;
assign t[328] = 6083;
assign s[329] = 14455085;
assign t[329] = 6078;
assign s[330] = 14449007;
assign t[330] = 6073;
assign s[331] = 14442933;
assign t[331] = 6068;
assign s[332] = 14436865;
assign t[332] = 6063;
assign s[333] = 14430801;
assign t[333] = 6058;
assign s[334] = 14424743;
assign t[334] = 6053;
assign s[335] = 14418690;
assign t[335] = 6048;
assign s[336] = 14412642;
assign t[336] = 6043;
assign s[337] = 14406599;
assign t[337] = 6037;
assign s[338] = 14400561;
assign t[338] = 6032;
assign s[339] = 14394528;
assign t[339] = 6027;
assign s[340] = 14388500;
assign t[340] = 6022;
assign s[341] = 14382477;
assign t[341] = 6017;
assign s[342] = 14376459;
assign t[342] = 6012;
assign s[343] = 14370447;
assign t[343] = 6007;
assign s[344] = 14364439;
assign t[344] = 6002;
assign s[345] = 14358436;
assign t[345] = 5997;
assign s[346] = 14352439;
assign t[346] = 5992;
assign s[347] = 14346446;
assign t[347] = 5987;
assign s[348] = 14340458;
assign t[348] = 5982;
assign s[349] = 14334476;
assign t[349] = 5977;
assign s[350] = 14328498;
assign t[350] = 5972;
assign s[351] = 14322525;
assign t[351] = 5967;
assign s[352] = 14316558;
assign t[352] = 5962;
assign s[353] = 14310595;
assign t[353] = 5957;
assign s[354] = 14304637;
assign t[354] = 5952;
assign s[355] = 14298684;
assign t[355] = 5947;
assign s[356] = 14292736;
assign t[356] = 5942;
assign s[357] = 14286793;
assign t[357] = 5937;
assign s[358] = 14280855;
assign t[358] = 5933;
assign s[359] = 14274922;
assign t[359] = 5928;
assign s[360] = 14268994;
assign t[360] = 5923;
assign s[361] = 14263071;
assign t[361] = 5918;
assign s[362] = 14257153;
assign t[362] = 5913;
assign s[363] = 14251239;
assign t[363] = 5908;
assign s[364] = 14245331;
assign t[364] = 5903;
assign s[365] = 14239427;
assign t[365] = 5898;
assign s[366] = 14233529;
assign t[366] = 5893;
assign s[367] = 14227635;
assign t[367] = 5888;
assign s[368] = 14221746;
assign t[368] = 5884;
assign s[369] = 14215862;
assign t[369] = 5879;
assign s[370] = 14209983;
assign t[370] = 5874;
assign s[371] = 14204108;
assign t[371] = 5869;
assign s[372] = 14198239;
assign t[372] = 5864;
assign s[373] = 14192374;
assign t[373] = 5859;
assign s[374] = 14186514;
assign t[374] = 5854;
assign s[375] = 14180660;
assign t[375] = 5850;
assign s[376] = 14174809;
assign t[376] = 5845;
assign s[377] = 14168964;
assign t[377] = 5840;
assign s[378] = 14163124;
assign t[378] = 5835;
assign s[379] = 14157288;
assign t[379] = 5830;
assign s[380] = 14151457;
assign t[380] = 5826;
assign s[381] = 14145631;
assign t[381] = 5821;
assign s[382] = 14139810;
assign t[382] = 5816;
assign s[383] = 14133993;
assign t[383] = 5811;
assign s[384] = 14128182;
assign t[384] = 5806;
assign s[385] = 14122375;
assign t[385] = 5802;
assign s[386] = 14116573;
assign t[386] = 5797;
assign s[387] = 14110775;
assign t[387] = 5792;
assign s[388] = 14104983;
assign t[388] = 5787;
assign s[389] = 14099195;
assign t[389] = 5783;
assign s[390] = 14093412;
assign t[390] = 5778;
assign s[391] = 14087634;
assign t[391] = 5773;
assign s[392] = 14081860;
assign t[392] = 5768;
assign s[393] = 14076091;
assign t[393] = 5764;
assign s[394] = 14070327;
assign t[394] = 5759;
assign s[395] = 14064567;
assign t[395] = 5754;
assign s[396] = 14058813;
assign t[396] = 5750;
assign s[397] = 14053063;
assign t[397] = 5745;
assign s[398] = 14047317;
assign t[398] = 5740;
assign s[399] = 14041577;
assign t[399] = 5735;
assign s[400] = 14035841;
assign t[400] = 5731;
assign s[401] = 14030109;
assign t[401] = 5726;
assign s[402] = 14024383;
assign t[402] = 5721;
assign s[403] = 14018661;
assign t[403] = 5717;
assign s[404] = 14012944;
assign t[404] = 5712;
assign s[405] = 14007231;
assign t[405] = 5707;
assign s[406] = 14001523;
assign t[406] = 5703;
assign s[407] = 13995820;
assign t[407] = 5698;
assign s[408] = 13990121;
assign t[408] = 5693;
assign s[409] = 13984427;
assign t[409] = 5689;
assign s[410] = 13978738;
assign t[410] = 5684;
assign s[411] = 13973053;
assign t[411] = 5680;
assign s[412] = 13967373;
assign t[412] = 5675;
assign s[413] = 13961698;
assign t[413] = 5670;
assign s[414] = 13956027;
assign t[414] = 5666;
assign s[415] = 13950361;
assign t[415] = 5661;
assign s[416] = 13944699;
assign t[416] = 5657;
assign s[417] = 13939042;
assign t[417] = 5652;
assign s[418] = 13933389;
assign t[418] = 5647;
assign s[419] = 13927741;
assign t[419] = 5643;
assign s[420] = 13922098;
assign t[420] = 5638;
assign s[421] = 13916459;
assign t[421] = 5634;
assign s[422] = 13910825;
assign t[422] = 5629;
assign s[423] = 13905196;
assign t[423] = 5625;
assign s[424] = 13899570;
assign t[424] = 5620;
assign s[425] = 13893950;
assign t[425] = 5615;
assign s[426] = 13888334;
assign t[426] = 5611;
assign s[427] = 13882723;
assign t[427] = 5606;
assign s[428] = 13877116;
assign t[428] = 5602;
assign s[429] = 13871513;
assign t[429] = 5597;
assign s[430] = 13865915;
assign t[430] = 5593;
assign s[431] = 13860322;
assign t[431] = 5588;
assign s[432] = 13854733;
assign t[432] = 5584;
assign s[433] = 13849149;
assign t[433] = 5579;
assign s[434] = 13843569;
assign t[434] = 5575;
assign s[435] = 13837994;
assign t[435] = 5570;
assign s[436] = 13832423;
assign t[436] = 5566;
assign s[437] = 13826856;
assign t[437] = 5561;
assign s[438] = 13821295;
assign t[438] = 5557;
assign s[439] = 13815737;
assign t[439] = 5552;
assign s[440] = 13810184;
assign t[440] = 5548;
assign s[441] = 13804636;
assign t[441] = 5544;
assign s[442] = 13799092;
assign t[442] = 5539;
assign s[443] = 13793552;
assign t[443] = 5535;
assign s[444] = 13788017;
assign t[444] = 5530;
assign s[445] = 13782486;
assign t[445] = 5526;
assign s[446] = 13776960;
assign t[446] = 5521;
assign s[447] = 13771438;
assign t[447] = 5517;
assign s[448] = 13765921;
assign t[448] = 5512;
assign s[449] = 13760408;
assign t[449] = 5508;
assign s[450] = 13754899;
assign t[450] = 5504;
assign s[451] = 13749395;
assign t[451] = 5499;
assign s[452] = 13743895;
assign t[452] = 5495;
assign s[453] = 13738400;
assign t[453] = 5490;
assign s[454] = 13732909;
assign t[454] = 5486;
assign s[455] = 13727422;
assign t[455] = 5482;
assign s[456] = 13721940;
assign t[456] = 5477;
assign s[457] = 13716462;
assign t[457] = 5473;
assign s[458] = 13710989;
assign t[458] = 5469;
assign s[459] = 13705520;
assign t[459] = 5464;
assign s[460] = 13700055;
assign t[460] = 5460;
assign s[461] = 13694595;
assign t[461] = 5456;
assign s[462] = 13689139;
assign t[462] = 5451;
assign s[463] = 13683687;
assign t[463] = 5447;
assign s[464] = 13678240;
assign t[464] = 5442;
assign s[465] = 13672797;
assign t[465] = 5438;
assign s[466] = 13667358;
assign t[466] = 5434;
assign s[467] = 13661924;
assign t[467] = 5430;
assign s[468] = 13656494;
assign t[468] = 5425;
assign s[469] = 13651068;
assign t[469] = 5421;
assign s[470] = 13645647;
assign t[470] = 5417;
assign s[471] = 13640230;
assign t[471] = 5412;
assign s[472] = 13634817;
assign t[472] = 5408;
assign s[473] = 13629408;
assign t[473] = 5404;
assign s[474] = 13624004;
assign t[474] = 5399;
assign s[475] = 13618604;
assign t[475] = 5395;
assign s[476] = 13613209;
assign t[476] = 5391;
assign s[477] = 13607817;
assign t[477] = 5387;
assign s[478] = 13602430;
assign t[478] = 5382;
assign s[479] = 13597047;
assign t[479] = 5378;
assign s[480] = 13591669;
assign t[480] = 5374;
assign s[481] = 13586294;
assign t[481] = 5370;
assign s[482] = 13580924;
assign t[482] = 5365;
assign s[483] = 13575558;
assign t[483] = 5361;
assign s[484] = 13570197;
assign t[484] = 5357;
assign s[485] = 13564839;
assign t[485] = 5353;
assign s[486] = 13559486;
assign t[486] = 5348;
assign s[487] = 13554137;
assign t[487] = 5344;
assign s[488] = 13548793;
assign t[488] = 5340;
assign s[489] = 13543452;
assign t[489] = 5336;
assign s[490] = 13538116;
assign t[490] = 5332;
assign s[491] = 13532784;
assign t[491] = 5327;
assign s[492] = 13527456;
assign t[492] = 5323;
assign s[493] = 13522132;
assign t[493] = 5319;
assign s[494] = 13516813;
assign t[494] = 5315;
assign s[495] = 13511498;
assign t[495] = 5311;
assign s[496] = 13506186;
assign t[496] = 5306;
assign s[497] = 13500879;
assign t[497] = 5302;
assign s[498] = 13495577;
assign t[498] = 5298;
assign s[499] = 13490278;
assign t[499] = 5294;
assign s[500] = 13484984;
assign t[500] = 5290;
assign s[501] = 13479693;
assign t[501] = 5286;
assign s[502] = 13474407;
assign t[502] = 5282;
assign s[503] = 13469125;
assign t[503] = 5277;
assign s[504] = 13463847;
assign t[504] = 5273;
assign s[505] = 13458574;
assign t[505] = 5269;
assign s[506] = 13453304;
assign t[506] = 5265;
assign s[507] = 13448038;
assign t[507] = 5261;
assign s[508] = 13442777;
assign t[508] = 5257;
assign s[509] = 13437520;
assign t[509] = 5253;
assign s[510] = 13432267;
assign t[510] = 5249;
assign s[511] = 13427018;
assign t[511] = 5244;
assign s[512] = 13421773;
assign t[512] = 5240;
assign s[513] = 13416532;
assign t[513] = 5236;
assign s[514] = 13411295;
assign t[514] = 5232;
assign s[515] = 13406063;
assign t[515] = 5228;
assign s[516] = 13400834;
assign t[516] = 5224;
assign s[517] = 13395609;
assign t[517] = 5220;
assign s[518] = 13390389;
assign t[518] = 5216;
assign s[519] = 13385173;
assign t[519] = 5212;
assign s[520] = 13379960;
assign t[520] = 5208;
assign s[521] = 13374752;
assign t[521] = 5204;
assign s[522] = 13369548;
assign t[522] = 5200;
assign s[523] = 13364348;
assign t[523] = 5196;
assign s[524] = 13359152;
assign t[524] = 5192;
assign s[525] = 13353960;
assign t[525] = 5188;
assign s[526] = 13348772;
assign t[526] = 5183;
assign s[527] = 13343588;
assign t[527] = 5179;
assign s[528] = 13338408;
assign t[528] = 5175;
assign s[529] = 13333232;
assign t[529] = 5171;
assign s[530] = 13328060;
assign t[530] = 5167;
assign s[531] = 13322892;
assign t[531] = 5163;
assign s[532] = 13317728;
assign t[532] = 5159;
assign s[533] = 13312568;
assign t[533] = 5155;
assign s[534] = 13307412;
assign t[534] = 5151;
assign s[535] = 13302260;
assign t[535] = 5147;
assign s[536] = 13297112;
assign t[536] = 5143;
assign s[537] = 13291968;
assign t[537] = 5139;
assign s[538] = 13286828;
assign t[538] = 5135;
assign s[539] = 13281692;
assign t[539] = 5132;
assign s[540] = 13276560;
assign t[540] = 5128;
assign s[541] = 13271432;
assign t[541] = 5124;
assign s[542] = 13266308;
assign t[542] = 5120;
assign s[543] = 13261188;
assign t[543] = 5116;
assign s[544] = 13256072;
assign t[544] = 5112;
assign s[545] = 13250960;
assign t[545] = 5108;
assign s[546] = 13245851;
assign t[546] = 5104;
assign s[547] = 13240747;
assign t[547] = 5100;
assign s[548] = 13235647;
assign t[548] = 5096;
assign s[549] = 13230550;
assign t[549] = 5092;
assign s[550] = 13225457;
assign t[550] = 5088;
assign s[551] = 13220369;
assign t[551] = 5084;
assign s[552] = 13215284;
assign t[552] = 5080;
assign s[553] = 13210203;
assign t[553] = 5076;
assign s[554] = 13205126;
assign t[554] = 5073;
assign s[555] = 13200053;
assign t[555] = 5069;
assign s[556] = 13194984;
assign t[556] = 5065;
assign s[557] = 13189919;
assign t[557] = 5061;
assign s[558] = 13184857;
assign t[558] = 5057;
assign s[559] = 13179800;
assign t[559] = 5053;
assign s[560] = 13174746;
assign t[560] = 5049;
assign s[561] = 13169697;
assign t[561] = 5045;
assign s[562] = 13164651;
assign t[562] = 5041;
assign s[563] = 13159609;
assign t[563] = 5038;
assign s[564] = 13154571;
assign t[564] = 5034;
assign s[565] = 13149536;
assign t[565] = 5030;
assign s[566] = 13144506;
assign t[566] = 5026;
assign s[567] = 13139479;
assign t[567] = 5022;
assign s[568] = 13134457;
assign t[568] = 5018;
assign s[569] = 13129438;
assign t[569] = 5015;
assign s[570] = 13124423;
assign t[570] = 5011;
assign s[571] = 13119411;
assign t[571] = 5007;
assign s[572] = 13114404;
assign t[572] = 5003;
assign s[573] = 13109400;
assign t[573] = 4999;
assign s[574] = 13104401;
assign t[574] = 4995;
assign s[575] = 13099405;
assign t[575] = 4992;
assign s[576] = 13094413;
assign t[576] = 4988;
assign s[577] = 13089424;
assign t[577] = 4984;
assign s[578] = 13084440;
assign t[578] = 4980;
assign s[579] = 13079459;
assign t[579] = 4976;
assign s[580] = 13074482;
assign t[580] = 4973;
assign s[581] = 13069509;
assign t[581] = 4969;
assign s[582] = 13064539;
assign t[582] = 4965;
assign s[583] = 13059574;
assign t[583] = 4961;
assign s[584] = 13054612;
assign t[584] = 4958;
assign s[585] = 13049654;
assign t[585] = 4954;
assign s[586] = 13044699;
assign t[586] = 4950;
assign s[587] = 13039749;
assign t[587] = 4946;
assign s[588] = 13034802;
assign t[588] = 4943;
assign s[589] = 13029859;
assign t[589] = 4939;
assign s[590] = 13024920;
assign t[590] = 4935;
assign s[591] = 13019984;
assign t[591] = 4931;
assign s[592] = 13015052;
assign t[592] = 4928;
assign s[593] = 13010124;
assign t[593] = 4924;
assign s[594] = 13005200;
assign t[594] = 4920;
assign s[595] = 13000279;
assign t[595] = 4916;
assign s[596] = 12995363;
assign t[596] = 4913;
assign s[597] = 12990449;
assign t[597] = 4909;
assign s[598] = 12985540;
assign t[598] = 4905;
assign s[599] = 12980634;
assign t[599] = 4902;
assign s[600] = 12975732;
assign t[600] = 4898;
assign s[601] = 12970834;
assign t[601] = 4894;
assign s[602] = 12965939;
assign t[602] = 4890;
assign s[603] = 12961048;
assign t[603] = 4887;
assign s[604] = 12956161;
assign t[604] = 4883;
assign s[605] = 12951277;
assign t[605] = 4879;
assign s[606] = 12946397;
assign t[606] = 4876;
assign s[607] = 12941521;
assign t[607] = 4872;
assign s[608] = 12936649;
assign t[608] = 4868;
assign s[609] = 12931780;
assign t[609] = 4865;
assign s[610] = 12926914;
assign t[610] = 4861;
assign s[611] = 12922053;
assign t[611] = 4857;
assign s[612] = 12917195;
assign t[612] = 4854;
assign s[613] = 12912341;
assign t[613] = 4850;
assign s[614] = 12907490;
assign t[614] = 4846;
assign s[615] = 12902643;
assign t[615] = 4843;
assign s[616] = 12897800;
assign t[616] = 4839;
assign s[617] = 12892960;
assign t[617] = 4836;
assign s[618] = 12888124;
assign t[618] = 4832;
assign s[619] = 12883292;
assign t[619] = 4828;
assign s[620] = 12878463;
assign t[620] = 4825;
assign s[621] = 12873638;
assign t[621] = 4821;
assign s[622] = 12868816;
assign t[622] = 4817;
assign s[623] = 12863998;
assign t[623] = 4814;
assign s[624] = 12859184;
assign t[624] = 4810;
assign s[625] = 12854373;
assign t[625] = 4807;
assign s[626] = 12849566;
assign t[626] = 4803;
assign s[627] = 12844762;
assign t[627] = 4799;
assign s[628] = 12839962;
assign t[628] = 4796;
assign s[629] = 12835166;
assign t[629] = 4792;
assign s[630] = 12830373;
assign t[630] = 4789;
assign s[631] = 12825584;
assign t[631] = 4785;
assign s[632] = 12820798;
assign t[632] = 4782;
assign s[633] = 12816016;
assign t[633] = 4778;
assign s[634] = 12811237;
assign t[634] = 4774;
assign s[635] = 12806462;
assign t[635] = 4771;
assign s[636] = 12801691;
assign t[636] = 4767;
assign s[637] = 12796923;
assign t[637] = 4764;
assign s[638] = 12792159;
assign t[638] = 4760;
assign s[639] = 12787398;
assign t[639] = 4757;
assign s[640] = 12782641;
assign t[640] = 4753;
assign s[641] = 12777887;
assign t[641] = 4750;
assign s[642] = 12773137;
assign t[642] = 4746;
assign s[643] = 12768390;
assign t[643] = 4743;
assign s[644] = 12763647;
assign t[644] = 4739;
assign s[645] = 12758908;
assign t[645] = 4736;
assign s[646] = 12754172;
assign t[646] = 4732;
assign s[647] = 12749439;
assign t[647] = 4729;
assign s[648] = 12744710;
assign t[648] = 4725;
assign s[649] = 12739985;
assign t[649] = 4722;
assign s[650] = 12735263;
assign t[650] = 4718;
assign s[651] = 12730544;
assign t[651] = 4715;
assign s[652] = 12725829;
assign t[652] = 4711;
assign s[653] = 12721118;
assign t[653] = 4708;
assign s[654] = 12716410;
assign t[654] = 4704;
assign s[655] = 12711705;
assign t[655] = 4701;
assign s[656] = 12707004;
assign t[656] = 4697;
assign s[657] = 12702306;
assign t[657] = 4694;
assign s[658] = 12697612;
assign t[658] = 4690;
assign s[659] = 12692922;
assign t[659] = 4687;
assign s[660] = 12688234;
assign t[660] = 4683;
assign s[661] = 12683551;
assign t[661] = 4680;
assign s[662] = 12678870;
assign t[662] = 4676;
assign s[663] = 12674193;
assign t[663] = 4673;
assign s[664] = 12669520;
assign t[664] = 4669;
assign s[665] = 12664850;
assign t[665] = 4666;
assign s[666] = 12660184;
assign t[666] = 4663;
assign s[667] = 12655521;
assign t[667] = 4659;
assign s[668] = 12650861;
assign t[668] = 4656;
assign s[669] = 12646205;
assign t[669] = 4652;
assign s[670] = 12641552;
assign t[670] = 4649;
assign s[671] = 12636903;
assign t[671] = 4645;
assign s[672] = 12632257;
assign t[672] = 4642;
assign s[673] = 12627614;
assign t[673] = 4639;
assign s[674] = 12622975;
assign t[674] = 4635;
assign s[675] = 12618340;
assign t[675] = 4632;
assign s[676] = 12613707;
assign t[676] = 4628;
assign s[677] = 12609078;
assign t[677] = 4625;
assign s[678] = 12604453;
assign t[678] = 4622;
assign s[679] = 12599831;
assign t[679] = 4618;
assign s[680] = 12595212;
assign t[680] = 4615;
assign s[681] = 12590597;
assign t[681] = 4611;
assign s[682] = 12585985;
assign t[682] = 4608;
assign s[683] = 12581376;
assign t[683] = 4605;
assign s[684] = 12576771;
assign t[684] = 4601;
assign s[685] = 12572169;
assign t[685] = 4598;
assign s[686] = 12567571;
assign t[686] = 4595;
assign s[687] = 12562976;
assign t[687] = 4591;
assign s[688] = 12558384;
assign t[688] = 4588;
assign s[689] = 12553796;
assign t[689] = 4585;
assign s[690] = 12549211;
assign t[690] = 4581;
assign s[691] = 12544629;
assign t[691] = 4578;
assign s[692] = 12540051;
assign t[692] = 4574;
assign s[693] = 12535476;
assign t[693] = 4571;
assign s[694] = 12530904;
assign t[694] = 4568;
assign s[695] = 12526336;
assign t[695] = 4564;
assign s[696] = 12521771;
assign t[696] = 4561;
assign s[697] = 12517209;
assign t[697] = 4558;
assign s[698] = 12512651;
assign t[698] = 4555;
assign s[699] = 12508096;
assign t[699] = 4551;
assign s[700] = 12503544;
assign t[700] = 4548;
assign s[701] = 12498995;
assign t[701] = 4545;
assign s[702] = 12494450;
assign t[702] = 4541;
assign s[703] = 12489909;
assign t[703] = 4538;
assign s[704] = 12485370;
assign t[704] = 4535;
assign s[705] = 12480835;
assign t[705] = 4531;
assign s[706] = 12476303;
assign t[706] = 4528;
assign s[707] = 12471774;
assign t[707] = 4525;
assign s[708] = 12467249;
assign t[708] = 4522;
assign s[709] = 12462727;
assign t[709] = 4518;
assign s[710] = 12458208;
assign t[710] = 4515;
assign s[711] = 12453693;
assign t[711] = 4512;
assign s[712] = 12449181;
assign t[712] = 4508;
assign s[713] = 12444672;
assign t[713] = 4505;
assign s[714] = 12440166;
assign t[714] = 4502;
assign s[715] = 12435664;
assign t[715] = 4499;
assign s[716] = 12431164;
assign t[716] = 4495;
assign s[717] = 12426669;
assign t[717] = 4492;
assign s[718] = 12422176;
assign t[718] = 4489;
assign s[719] = 12417687;
assign t[719] = 4486;
assign s[720] = 12413200;
assign t[720] = 4482;
assign s[721] = 12408717;
assign t[721] = 4479;
assign s[722] = 12404238;
assign t[722] = 4476;
assign s[723] = 12399761;
assign t[723] = 4473;
assign s[724] = 12395288;
assign t[724] = 4469;
assign s[725] = 12390818;
assign t[725] = 4466;
assign s[726] = 12386351;
assign t[726] = 4463;
assign s[727] = 12381888;
assign t[727] = 4460;
assign s[728] = 12377427;
assign t[728] = 4457;
assign s[729] = 12372970;
assign t[729] = 4453;
assign s[730] = 12368516;
assign t[730] = 4450;
assign s[731] = 12364066;
assign t[731] = 4447;
assign s[732] = 12359618;
assign t[732] = 4444;
assign s[733] = 12355174;
assign t[733] = 4441;
assign s[734] = 12350733;
assign t[734] = 4437;
assign s[735] = 12346295;
assign t[735] = 4434;
assign s[736] = 12341860;
assign t[736] = 4431;
assign s[737] = 12337429;
assign t[737] = 4428;
assign s[738] = 12333000;
assign t[738] = 4425;
assign s[739] = 12328575;
assign t[739] = 4422;
assign s[740] = 12324153;
assign t[740] = 4418;
assign s[741] = 12319734;
assign t[741] = 4415;
assign s[742] = 12315319;
assign t[742] = 4412;
assign s[743] = 12310906;
assign t[743] = 4409;
assign s[744] = 12306497;
assign t[744] = 4406;
assign s[745] = 12302090;
assign t[745] = 4403;
assign s[746] = 12297687;
assign t[746] = 4399;
assign s[747] = 12293288;
assign t[747] = 4396;
assign s[748] = 12288891;
assign t[748] = 4393;
assign s[749] = 12284497;
assign t[749] = 4390;
assign s[750] = 12280107;
assign t[750] = 4387;
assign s[751] = 12275719;
assign t[751] = 4384;
assign s[752] = 12271335;
assign t[752] = 4381;
assign s[753] = 12266954;
assign t[753] = 4377;
assign s[754] = 12262576;
assign t[754] = 4374;
assign s[755] = 12258201;
assign t[755] = 4371;
assign s[756] = 12253830;
assign t[756] = 4368;
assign s[757] = 12249461;
assign t[757] = 4365;
assign s[758] = 12245096;
assign t[758] = 4362;
assign s[759] = 12240733;
assign t[759] = 4359;
assign s[760] = 12236374;
assign t[760] = 4356;
assign s[761] = 12232018;
assign t[761] = 4353;
assign s[762] = 12227665;
assign t[762] = 4349;
assign s[763] = 12223315;
assign t[763] = 4346;
assign s[764] = 12218968;
assign t[764] = 4343;
assign s[765] = 12214624;
assign t[765] = 4340;
assign s[766] = 12210284;
assign t[766] = 4337;
assign s[767] = 12205946;
assign t[767] = 4334;
assign s[768] = 12201612;
assign t[768] = 4331;
assign s[769] = 12197280;
assign t[769] = 4328;
assign s[770] = 12192952;
assign t[770] = 4325;
assign s[771] = 12188627;
assign t[771] = 4322;
assign s[772] = 12184305;
assign t[772] = 4319;
assign s[773] = 12179985;
assign t[773] = 4316;
assign s[774] = 12175669;
assign t[774] = 4313;
assign s[775] = 12171356;
assign t[775] = 4309;
assign s[776] = 12167046;
assign t[776] = 4306;
assign s[777] = 12162739;
assign t[777] = 4303;
assign s[778] = 12158435;
assign t[778] = 4300;
assign s[779] = 12154135;
assign t[779] = 4297;
assign s[780] = 12149837;
assign t[780] = 4294;
assign s[781] = 12145542;
assign t[781] = 4291;
assign s[782] = 12141250;
assign t[782] = 4288;
assign s[783] = 12136962;
assign t[783] = 4285;
assign s[784] = 12132676;
assign t[784] = 4282;
assign s[785] = 12128393;
assign t[785] = 4279;
assign s[786] = 12124114;
assign t[786] = 4276;
assign s[787] = 12119837;
assign t[787] = 4273;
assign s[788] = 12115564;
assign t[788] = 4270;
assign s[789] = 12111293;
assign t[789] = 4267;
assign s[790] = 12107026;
assign t[790] = 4264;
assign s[791] = 12102761;
assign t[791] = 4261;
assign s[792] = 12098500;
assign t[792] = 4258;
assign s[793] = 12094241;
assign t[793] = 4255;
assign s[794] = 12089985;
assign t[794] = 4252;
assign s[795] = 12085733;
assign t[795] = 4249;
assign s[796] = 12081483;
assign t[796] = 4246;
assign s[797] = 12077237;
assign t[797] = 4243;
assign s[798] = 12072993;
assign t[798] = 4240;
assign s[799] = 12068753;
assign t[799] = 4237;
assign s[800] = 12064515;
assign t[800] = 4234;
assign s[801] = 12060280;
assign t[801] = 4231;
assign s[802] = 12056049;
assign t[802] = 4228;
assign s[803] = 12051820;
assign t[803] = 4225;
assign s[804] = 12047594;
assign t[804] = 4222;
assign s[805] = 12043371;
assign t[805] = 4219;
assign s[806] = 12039152;
assign t[806] = 4216;
assign s[807] = 12034935;
assign t[807] = 4213;
assign s[808] = 12030721;
assign t[808] = 4210;
assign s[809] = 12026510;
assign t[809] = 4208;
assign s[810] = 12022302;
assign t[810] = 4205;
assign s[811] = 12018097;
assign t[811] = 4202;
assign s[812] = 12013895;
assign t[812] = 4199;
assign s[813] = 12009695;
assign t[813] = 4196;
assign s[814] = 12005499;
assign t[814] = 4193;
assign s[815] = 12001306;
assign t[815] = 4190;
assign s[816] = 11997115;
assign t[816] = 4187;
assign s[817] = 11992928;
assign t[817] = 4184;
assign s[818] = 11988743;
assign t[818] = 4181;
assign s[819] = 11984562;
assign t[819] = 4178;
assign s[820] = 11980383;
assign t[820] = 4175;
assign s[821] = 11976207;
assign t[821] = 4172;
assign s[822] = 11972034;
assign t[822] = 4169;
assign s[823] = 11967864;
assign t[823] = 4167;
assign s[824] = 11963697;
assign t[824] = 4164;
assign s[825] = 11959533;
assign t[825] = 4161;
assign s[826] = 11955372;
assign t[826] = 4158;
assign s[827] = 11951213;
assign t[827] = 4155;
assign s[828] = 11947058;
assign t[828] = 4152;
assign s[829] = 11942905;
assign t[829] = 4149;
assign s[830] = 11938756;
assign t[830] = 4146;
assign s[831] = 11934609;
assign t[831] = 4143;
assign s[832] = 11930465;
assign t[832] = 4141;
assign s[833] = 11926324;
assign t[833] = 4138;
assign s[834] = 11922186;
assign t[834] = 4135;
assign s[835] = 11918050;
assign t[835] = 4132;
assign s[836] = 11913918;
assign t[836] = 4129;
assign s[837] = 11909788;
assign t[837] = 4126;
assign s[838] = 11905661;
assign t[838] = 4123;
assign s[839] = 11901538;
assign t[839] = 4121;
assign s[840] = 11897416;
assign t[840] = 4118;
assign s[841] = 11893298;
assign t[841] = 4115;
assign s[842] = 11889183;
assign t[842] = 4112;
assign s[843] = 11885070;
assign t[843] = 4109;
assign s[844] = 11880961;
assign t[844] = 4106;
assign s[845] = 11876854;
assign t[845] = 4103;
assign s[846] = 11872750;
assign t[846] = 4101;
assign s[847] = 11868649;
assign t[847] = 4098;
assign s[848] = 11864551;
assign t[848] = 4095;
assign s[849] = 11860455;
assign t[849] = 4092;
assign s[850] = 11856363;
assign t[850] = 4089;
assign s[851] = 11852273;
assign t[851] = 4086;
assign s[852] = 11848186;
assign t[852] = 4084;
assign s[853] = 11844102;
assign t[853] = 4081;
assign s[854] = 11840020;
assign t[854] = 4078;
assign s[855] = 11835942;
assign t[855] = 4075;
assign s[856] = 11831866;
assign t[856] = 4072;
assign s[857] = 11827793;
assign t[857] = 4070;
assign s[858] = 11823723;
assign t[858] = 4067;
assign s[859] = 11819656;
assign t[859] = 4064;
assign s[860] = 11815591;
assign t[860] = 4061;
assign s[861] = 11811529;
assign t[861] = 4058;
assign s[862] = 11807470;
assign t[862] = 4056;
assign s[863] = 11803414;
assign t[863] = 4053;
assign s[864] = 11799361;
assign t[864] = 4050;
assign s[865] = 11795310;
assign t[865] = 4047;
assign s[866] = 11791262;
assign t[866] = 4045;
assign s[867] = 11787217;
assign t[867] = 4042;
assign s[868] = 11783175;
assign t[868] = 4039;
assign s[869] = 11779136;
assign t[869] = 4036;
assign s[870] = 11775099;
assign t[870] = 4033;
assign s[871] = 11771065;
assign t[871] = 4031;
assign s[872] = 11767034;
assign t[872] = 4028;
assign s[873] = 11763005;
assign t[873] = 4025;
assign s[874] = 11758980;
assign t[874] = 4022;
assign s[875] = 11754957;
assign t[875] = 4020;
assign s[876] = 11750937;
assign t[876] = 4017;
assign s[877] = 11746919;
assign t[877] = 4014;
assign s[878] = 11742905;
assign t[878] = 4011;
assign s[879] = 11738893;
assign t[879] = 4009;
assign s[880] = 11734883;
assign t[880] = 4006;
assign s[881] = 11730877;
assign t[881] = 4003;
assign s[882] = 11726873;
assign t[882] = 4000;
assign s[883] = 11722872;
assign t[883] = 3998;
assign s[884] = 11718874;
assign t[884] = 3995;
assign s[885] = 11714879;
assign t[885] = 3992;
assign s[886] = 11710886;
assign t[886] = 3990;
assign s[887] = 11706896;
assign t[887] = 3987;
assign s[888] = 11702908;
assign t[888] = 3984;
assign s[889] = 11698924;
assign t[889] = 3981;
assign s[890] = 11694942;
assign t[890] = 3979;
assign s[891] = 11690963;
assign t[891] = 3976;
assign s[892] = 11686986;
assign t[892] = 3973;
assign s[893] = 11683012;
assign t[893] = 3971;
assign s[894] = 11679041;
assign t[894] = 3968;
assign s[895] = 11675073;
assign t[895] = 3965;
assign s[896] = 11671107;
assign t[896] = 3963;
assign s[897] = 11667144;
assign t[897] = 3960;
assign s[898] = 11663184;
assign t[898] = 3957;
assign s[899] = 11659226;
assign t[899] = 3954;
assign s[900] = 11655271;
assign t[900] = 3952;
assign s[901] = 11651319;
assign t[901] = 3949;
assign s[902] = 11647369;
assign t[902] = 3946;
assign s[903] = 11643422;
assign t[903] = 3944;
assign s[904] = 11639478;
assign t[904] = 3941;
assign s[905] = 11635536;
assign t[905] = 3938;
assign s[906] = 11631597;
assign t[906] = 3936;
assign s[907] = 11627661;
assign t[907] = 3933;
assign s[908] = 11623728;
assign t[908] = 3930;
assign s[909] = 11619797;
assign t[909] = 3928;
assign s[910] = 11615868;
assign t[910] = 3925;
assign s[911] = 11611943;
assign t[911] = 3922;
assign s[912] = 11608020;
assign t[912] = 3920;
assign s[913] = 11604100;
assign t[913] = 3917;
assign s[914] = 11600182;
assign t[914] = 3915;
assign s[915] = 11596267;
assign t[915] = 3912;
assign s[916] = 11592355;
assign t[916] = 3909;
assign s[917] = 11588445;
assign t[917] = 3907;
assign s[918] = 11584538;
assign t[918] = 3904;
assign s[919] = 11580633;
assign t[919] = 3901;
assign s[920] = 11576731;
assign t[920] = 3899;
assign s[921] = 11572832;
assign t[921] = 3896;
assign s[922] = 11568936;
assign t[922] = 3893;
assign s[923] = 11565042;
assign t[923] = 3891;
assign s[924] = 11561150;
assign t[924] = 3888;
assign s[925] = 11557262;
assign t[925] = 3886;
assign s[926] = 11553376;
assign t[926] = 3883;
assign s[927] = 11549492;
assign t[927] = 3880;
assign s[928] = 11545611;
assign t[928] = 3878;
assign s[929] = 11541733;
assign t[929] = 3875;
assign s[930] = 11537857;
assign t[930] = 3873;
assign s[931] = 11533984;
assign t[931] = 3870;
assign s[932] = 11530114;
assign t[932] = 3867;
assign s[933] = 11526246;
assign t[933] = 3865;
assign s[934] = 11522381;
assign t[934] = 3862;
assign s[935] = 11518518;
assign t[935] = 3860;
assign s[936] = 11514658;
assign t[936] = 3857;
assign s[937] = 11510800;
assign t[937] = 3854;
assign s[938] = 11506945;
assign t[938] = 3852;
assign s[939] = 11503093;
assign t[939] = 3849;
assign s[940] = 11499243;
assign t[940] = 3847;
assign s[941] = 11495396;
assign t[941] = 3844;
assign s[942] = 11491551;
assign t[942] = 3842;
assign s[943] = 11487709;
assign t[943] = 3839;
assign s[944] = 11483870;
assign t[944] = 3836;
assign s[945] = 11480033;
assign t[945] = 3834;
assign s[946] = 11476199;
assign t[946] = 3831;
assign s[947] = 11472367;
assign t[947] = 3829;
assign s[948] = 11468538;
assign t[948] = 3826;
assign s[949] = 11464711;
assign t[949] = 3824;
assign s[950] = 11460887;
assign t[950] = 3821;
assign s[951] = 11457065;
assign t[951] = 3819;
assign s[952] = 11453246;
assign t[952] = 3816;
assign s[953] = 11449430;
assign t[953] = 3813;
assign s[954] = 11445616;
assign t[954] = 3811;
assign s[955] = 11441805;
assign t[955] = 3808;
assign s[956] = 11437996;
assign t[956] = 3806;
assign s[957] = 11434189;
assign t[957] = 3803;
assign s[958] = 11430386;
assign t[958] = 3801;
assign s[959] = 11426584;
assign t[959] = 3798;
assign s[960] = 11422786;
assign t[960] = 3796;
assign s[961] = 11418989;
assign t[961] = 3793;
assign s[962] = 11415196;
assign t[962] = 3791;
assign s[963] = 11411404;
assign t[963] = 3788;
assign s[964] = 11407616;
assign t[964] = 3786;
assign s[965] = 11403830;
assign t[965] = 3783;
assign s[966] = 11400046;
assign t[966] = 3781;
assign s[967] = 11396265;
assign t[967] = 3778;
assign s[968] = 11392486;
assign t[968] = 3776;
assign s[969] = 11388710;
assign t[969] = 3773;
assign s[970] = 11384937;
assign t[970] = 3771;
assign s[971] = 11381166;
assign t[971] = 3768;
assign s[972] = 11377397;
assign t[972] = 3766;
assign s[973] = 11373631;
assign t[973] = 3763;
assign s[974] = 11369867;
assign t[974] = 3761;
assign s[975] = 11366106;
assign t[975] = 3758;
assign s[976] = 11362348;
assign t[976] = 3756;
assign s[977] = 11358591;
assign t[977] = 3753;
assign s[978] = 11354838;
assign t[978] = 3751;
assign s[979] = 11351087;
assign t[979] = 3748;
assign s[980] = 11347338;
assign t[980] = 3746;
assign s[981] = 11343592;
assign t[981] = 3743;
assign s[982] = 11339848;
assign t[982] = 3741;
assign s[983] = 11336107;
assign t[983] = 3738;
assign s[984] = 11332368;
assign t[984] = 3736;
assign s[985] = 11328631;
assign t[985] = 3733;
assign s[986] = 11324897;
assign t[986] = 3731;
assign s[987] = 11321166;
assign t[987] = 3728;
assign s[988] = 11317437;
assign t[988] = 3726;
assign s[989] = 11313711;
assign t[989] = 3724;
assign s[990] = 11309986;
assign t[990] = 3721;
assign s[991] = 11306265;
assign t[991] = 3719;
assign s[992] = 11302546;
assign t[992] = 3716;
assign s[993] = 11298829;
assign t[993] = 3714;
assign s[994] = 11295115;
assign t[994] = 3711;
assign s[995] = 11291403;
assign t[995] = 3709;
assign s[996] = 11287693;
assign t[996] = 3706;
assign s[997] = 11283987;
assign t[997] = 3704;
assign s[998] = 11280282;
assign t[998] = 3702;
assign s[999] = 11276580;
assign t[999] = 3699;
assign s[1000] = 11272880;
assign t[1000] = 3697;
assign s[1001] = 11269183;
assign t[1001] = 3694;
assign s[1002] = 11265488;
assign t[1002] = 3692;
assign s[1003] = 11261796;
assign t[1003] = 3689;
assign s[1004] = 11258106;
assign t[1004] = 3687;
assign s[1005] = 11254418;
assign t[1005] = 3685;
assign s[1006] = 11250733;
assign t[1006] = 3682;
assign s[1007] = 11247050;
assign t[1007] = 3680;
assign s[1008] = 11243370;
assign t[1008] = 3677;
assign s[1009] = 11239692;
assign t[1009] = 3675;
assign s[1010] = 11236017;
assign t[1010] = 3673;
assign s[1011] = 11232344;
assign t[1011] = 3670;
assign s[1012] = 11228673;
assign t[1012] = 3668;
assign s[1013] = 11225005;
assign t[1013] = 3665;
assign s[1014] = 11221339;
assign t[1014] = 3663;
assign s[1015] = 11217675;
assign t[1015] = 3661;
assign s[1016] = 11214014;
assign t[1016] = 3658;
assign s[1017] = 11210355;
assign t[1017] = 3656;
assign s[1018] = 11206699;
assign t[1018] = 3653;
assign s[1019] = 11203045;
assign t[1019] = 3651;
assign s[1020] = 11199393;
assign t[1020] = 3649;
assign s[1021] = 11195744;
assign t[1021] = 3646;
assign s[1022] = 11192097;
assign t[1022] = 3644;
assign s[1023] = 11188453;
assign t[1023] = 3642;
assign s[1024] = 11184811;
assign t[1024] = 3639;
assign s[1025] = 11181171;
assign t[1025] = 3637;
assign s[1026] = 11177534;
assign t[1026] = 3634;
assign s[1027] = 11173899;
assign t[1027] = 3632;
assign s[1028] = 11170266;
assign t[1028] = 3630;
assign s[1029] = 11166636;
assign t[1029] = 3627;
assign s[1030] = 11163008;
assign t[1030] = 3625;
assign s[1031] = 11159383;
assign t[1031] = 3623;
assign s[1032] = 11155759;
assign t[1032] = 3620;
assign s[1033] = 11152139;
assign t[1033] = 3618;
assign s[1034] = 11148520;
assign t[1034] = 3616;
assign s[1035] = 11144904;
assign t[1035] = 3613;
assign s[1036] = 11141290;
assign t[1036] = 3611;
assign s[1037] = 11137679;
assign t[1037] = 3609;
assign s[1038] = 11134070;
assign t[1038] = 3606;
assign s[1039] = 11130463;
assign t[1039] = 3604;
assign s[1040] = 11126858;
assign t[1040] = 3602;
assign s[1041] = 11123256;
assign t[1041] = 3599;
assign s[1042] = 11119657;
assign t[1042] = 3597;
assign s[1043] = 11116059;
assign t[1043] = 3595;
assign s[1044] = 11112464;
assign t[1044] = 3592;
assign s[1045] = 11108871;
assign t[1045] = 3590;
assign s[1046] = 11105281;
assign t[1046] = 3588;
assign s[1047] = 11101693;
assign t[1047] = 3585;
assign s[1048] = 11098107;
assign t[1048] = 3583;
assign s[1049] = 11094523;
assign t[1049] = 3581;
assign s[1050] = 11090942;
assign t[1050] = 3578;
assign s[1051] = 11087363;
assign t[1051] = 3576;
assign s[1052] = 11083787;
assign t[1052] = 3574;
assign s[1053] = 11080213;
assign t[1053] = 3571;
assign s[1054] = 11076641;
assign t[1054] = 3569;
assign s[1055] = 11073071;
assign t[1055] = 3567;
assign s[1056] = 11069504;
assign t[1056] = 3565;
assign s[1057] = 11065938;
assign t[1057] = 3562;
assign s[1058] = 11062376;
assign t[1058] = 3560;
assign s[1059] = 11058815;
assign t[1059] = 3558;
assign s[1060] = 11055257;
assign t[1060] = 3555;
assign s[1061] = 11051701;
assign t[1061] = 3553;
assign s[1062] = 11048148;
assign t[1062] = 3551;
assign s[1063] = 11044596;
assign t[1063] = 3549;
assign s[1064] = 11041047;
assign t[1064] = 3546;
assign s[1065] = 11037500;
assign t[1065] = 3544;
assign s[1066] = 11033956;
assign t[1066] = 3542;
assign s[1067] = 11030414;
assign t[1067] = 3539;
assign s[1068] = 11026874;
assign t[1068] = 3537;
assign s[1069] = 11023336;
assign t[1069] = 3535;
assign s[1070] = 11019801;
assign t[1070] = 3533;
assign s[1071] = 11016268;
assign t[1071] = 3530;
assign s[1072] = 11012737;
assign t[1072] = 3528;
assign s[1073] = 11009208;
assign t[1073] = 3526;
assign s[1074] = 11005682;
assign t[1074] = 3524;
assign s[1075] = 11002158;
assign t[1075] = 3521;
assign s[1076] = 10998636;
assign t[1076] = 3519;
assign s[1077] = 10995116;
assign t[1077] = 3517;
assign s[1078] = 10991599;
assign t[1078] = 3515;
assign s[1079] = 10988084;
assign t[1079] = 3512;
assign s[1080] = 10984571;
assign t[1080] = 3510;
assign s[1081] = 10981061;
assign t[1081] = 3508;
assign s[1082] = 10977552;
assign t[1082] = 3506;
assign s[1083] = 10974046;
assign t[1083] = 3503;
assign s[1084] = 10970542;
assign t[1084] = 3501;
assign s[1085] = 10967041;
assign t[1085] = 3499;
assign s[1086] = 10963542;
assign t[1086] = 3497;
assign s[1087] = 10960044;
assign t[1087] = 3494;
assign s[1088] = 10956549;
assign t[1088] = 3492;
assign s[1089] = 10953057;
assign t[1089] = 3490;
assign s[1090] = 10949566;
assign t[1090] = 3488;
assign s[1091] = 10946078;
assign t[1091] = 3486;
assign s[1092] = 10942592;
assign t[1092] = 3483;
assign s[1093] = 10939108;
assign t[1093] = 3481;
assign s[1094] = 10935627;
assign t[1094] = 3479;
assign s[1095] = 10932147;
assign t[1095] = 3477;
assign s[1096] = 10928670;
assign t[1096] = 3474;
assign s[1097] = 10925195;
assign t[1097] = 3472;
assign s[1098] = 10921723;
assign t[1098] = 3470;
assign s[1099] = 10918252;
assign t[1099] = 3468;
assign s[1100] = 10914784;
assign t[1100] = 3466;
assign s[1101] = 10911318;
assign t[1101] = 3463;
assign s[1102] = 10907854;
assign t[1102] = 3461;
assign s[1103] = 10904392;
assign t[1103] = 3459;
assign s[1104] = 10900932;
assign t[1104] = 3457;
assign s[1105] = 10897475;
assign t[1105] = 3455;
assign s[1106] = 10894020;
assign t[1106] = 3452;
assign s[1107] = 10890567;
assign t[1107] = 3450;
assign s[1108] = 10887116;
assign t[1108] = 3448;
assign s[1109] = 10883668;
assign t[1109] = 3446;
assign s[1110] = 10880221;
assign t[1110] = 3444;
assign s[1111] = 10876777;
assign t[1111] = 3442;
assign s[1112] = 10873335;
assign t[1112] = 3439;
assign s[1113] = 10869895;
assign t[1113] = 3437;
assign s[1114] = 10866458;
assign t[1114] = 3435;
assign s[1115] = 10863022;
assign t[1115] = 3433;
assign s[1116] = 10859589;
assign t[1116] = 3431;
assign s[1117] = 10856158;
assign t[1117] = 3428;
assign s[1118] = 10852729;
assign t[1118] = 3426;
assign s[1119] = 10849302;
assign t[1119] = 3424;
assign s[1120] = 10845877;
assign t[1120] = 3422;
assign s[1121] = 10842455;
assign t[1121] = 3420;
assign s[1122] = 10839034;
assign t[1122] = 3418;
assign s[1123] = 10835616;
assign t[1123] = 3416;
assign s[1124] = 10832200;
assign t[1124] = 3413;
assign s[1125] = 10828786;
assign t[1125] = 3411;
assign s[1126] = 10825375;
assign t[1126] = 3409;
assign s[1127] = 10821965;
assign t[1127] = 3407;
assign s[1128] = 10818558;
assign t[1128] = 3405;
assign s[1129] = 10815152;
assign t[1129] = 3403;
assign s[1130] = 10811749;
assign t[1130] = 3400;
assign s[1131] = 10808348;
assign t[1131] = 3398;
assign s[1132] = 10804949;
assign t[1132] = 3396;
assign s[1133] = 10801553;
assign t[1133] = 3394;
assign s[1134] = 10798158;
assign t[1134] = 3392;
assign s[1135] = 10794766;
assign t[1135] = 3390;
assign s[1136] = 10791375;
assign t[1136] = 3388;
assign s[1137] = 10787987;
assign t[1137] = 3386;
assign s[1138] = 10784601;
assign t[1138] = 3383;
assign s[1139] = 10781217;
assign t[1139] = 3381;
assign s[1140] = 10777835;
assign t[1140] = 3379;
assign s[1141] = 10774456;
assign t[1141] = 3377;
assign s[1142] = 10771078;
assign t[1142] = 3375;
assign s[1143] = 10767703;
assign t[1143] = 3373;
assign s[1144] = 10764329;
assign t[1144] = 3371;
assign s[1145] = 10760958;
assign t[1145] = 3369;
assign s[1146] = 10757589;
assign t[1146] = 3367;
assign s[1147] = 10754222;
assign t[1147] = 3364;
assign s[1148] = 10750857;
assign t[1148] = 3362;
assign s[1149] = 10747494;
assign t[1149] = 3360;
assign s[1150] = 10744134;
assign t[1150] = 3358;
assign s[1151] = 10740775;
assign t[1151] = 3356;
assign s[1152] = 10737418;
assign t[1152] = 3354;
assign s[1153] = 10734064;
assign t[1153] = 3352;
assign s[1154] = 10730712;
assign t[1154] = 3350;
assign s[1155] = 10727362;
assign t[1155] = 3348;
assign s[1156] = 10724013;
assign t[1156] = 3346;
assign s[1157] = 10720667;
assign t[1157] = 3343;
assign s[1158] = 10717323;
assign t[1158] = 3341;
assign s[1159] = 10713982;
assign t[1159] = 3339;
assign s[1160] = 10710642;
assign t[1160] = 3337;
assign s[1161] = 10707304;
assign t[1161] = 3335;
assign s[1162] = 10703969;
assign t[1162] = 3333;
assign s[1163] = 10700635;
assign t[1163] = 3331;
assign s[1164] = 10697304;
assign t[1164] = 3329;
assign s[1165] = 10693974;
assign t[1165] = 3327;
assign s[1166] = 10690647;
assign t[1166] = 3325;
assign s[1167] = 10687322;
assign t[1167] = 3323;
assign s[1168] = 10683998;
assign t[1168] = 3321;
assign s[1169] = 10680677;
assign t[1169] = 3319;
assign s[1170] = 10677358;
assign t[1170] = 3316;
assign s[1171] = 10674041;
assign t[1171] = 3314;
assign s[1172] = 10670726;
assign t[1172] = 3312;
assign s[1173] = 10667414;
assign t[1173] = 3310;
assign s[1174] = 10664103;
assign t[1174] = 3308;
assign s[1175] = 10660794;
assign t[1175] = 3306;
assign s[1176] = 10657487;
assign t[1176] = 3304;
assign s[1177] = 10654183;
assign t[1177] = 3302;
assign s[1178] = 10650880;
assign t[1178] = 3300;
assign s[1179] = 10647580;
assign t[1179] = 3298;
assign s[1180] = 10644281;
assign t[1180] = 3296;
assign s[1181] = 10640985;
assign t[1181] = 3294;
assign s[1182] = 10637690;
assign t[1182] = 3292;
assign s[1183] = 10634398;
assign t[1183] = 3290;
assign s[1184] = 10631107;
assign t[1184] = 3288;
assign s[1185] = 10627819;
assign t[1185] = 3286;
assign s[1186] = 10624533;
assign t[1186] = 3284;
assign s[1187] = 10621249;
assign t[1187] = 3282;
assign s[1188] = 10617966;
assign t[1188] = 3280;
assign s[1189] = 10614686;
assign t[1189] = 3278;
assign s[1190] = 10611408;
assign t[1190] = 3276;
assign s[1191] = 10608132;
assign t[1191] = 3274;
assign s[1192] = 10604858;
assign t[1192] = 3272;
assign s[1193] = 10601586;
assign t[1193] = 3270;
assign s[1194] = 10598316;
assign t[1194] = 3268;
assign s[1195] = 10595048;
assign t[1195] = 3266;
assign s[1196] = 10591781;
assign t[1196] = 3264;
assign s[1197] = 10588517;
assign t[1197] = 3262;
assign s[1198] = 10585255;
assign t[1198] = 3260;
assign s[1199] = 10581995;
assign t[1199] = 3258;
assign s[1200] = 10578737;
assign t[1200] = 3255;
assign s[1201] = 10575481;
assign t[1201] = 3253;
assign s[1202] = 10572227;
assign t[1202] = 3251;
assign s[1203] = 10568975;
assign t[1203] = 3249;
assign s[1204] = 10565725;
assign t[1204] = 3247;
assign s[1205] = 10562477;
assign t[1205] = 3245;
assign s[1206] = 10559231;
assign t[1206] = 3244;
assign s[1207] = 10555987;
assign t[1207] = 3242;
assign s[1208] = 10552745;
assign t[1208] = 3240;
assign s[1209] = 10549505;
assign t[1209] = 3238;
assign s[1210] = 10546267;
assign t[1210] = 3236;
assign s[1211] = 10543031;
assign t[1211] = 3234;
assign s[1212] = 10539797;
assign t[1212] = 3232;
assign s[1213] = 10536565;
assign t[1213] = 3230;
assign s[1214] = 10533335;
assign t[1214] = 3228;
assign s[1215] = 10530107;
assign t[1215] = 3226;
assign s[1216] = 10526881;
assign t[1216] = 3224;
assign s[1217] = 10523657;
assign t[1217] = 3222;
assign s[1218] = 10520435;
assign t[1218] = 3220;
assign s[1219] = 10517214;
assign t[1219] = 3218;
assign s[1220] = 10513996;
assign t[1220] = 3216;
assign s[1221] = 10510780;
assign t[1221] = 3214;
assign s[1222] = 10507566;
assign t[1222] = 3212;
assign s[1223] = 10504353;
assign t[1223] = 3210;
assign s[1224] = 10501143;
assign t[1224] = 3208;
assign s[1225] = 10497934;
assign t[1225] = 3206;
assign s[1226] = 10494728;
assign t[1226] = 3204;
assign s[1227] = 10491523;
assign t[1227] = 3202;
assign s[1228] = 10488321;
assign t[1228] = 3200;
assign s[1229] = 10485120;
assign t[1229] = 3198;
assign s[1230] = 10481922;
assign t[1230] = 3196;
assign s[1231] = 10478725;
assign t[1231] = 3194;
assign s[1232] = 10475530;
assign t[1232] = 3192;
assign s[1233] = 10472337;
assign t[1233] = 3190;
assign s[1234] = 10469147;
assign t[1234] = 3188;
assign s[1235] = 10465958;
assign t[1235] = 3186;
assign s[1236] = 10462771;
assign t[1236] = 3185;
assign s[1237] = 10459586;
assign t[1237] = 3183;
assign s[1238] = 10456403;
assign t[1238] = 3181;
assign s[1239] = 10453222;
assign t[1239] = 3179;
assign s[1240] = 10450042;
assign t[1240] = 3177;
assign s[1241] = 10446865;
assign t[1241] = 3175;
assign s[1242] = 10443690;
assign t[1242] = 3173;
assign s[1243] = 10440516;
assign t[1243] = 3171;
assign s[1244] = 10437345;
assign t[1244] = 3169;
assign s[1245] = 10434175;
assign t[1245] = 3167;
assign s[1246] = 10431008;
assign t[1246] = 3165;
assign s[1247] = 10427842;
assign t[1247] = 3163;
assign s[1248] = 10424678;
assign t[1248] = 3161;
assign s[1249] = 10421516;
assign t[1249] = 3159;
assign s[1250] = 10418356;
assign t[1250] = 3158;
assign s[1251] = 10415198;
assign t[1251] = 3156;
assign s[1252] = 10412042;
assign t[1252] = 3154;
assign s[1253] = 10408888;
assign t[1253] = 3152;
assign s[1254] = 10405736;
assign t[1254] = 3150;
assign s[1255] = 10402585;
assign t[1255] = 3148;
assign s[1256] = 10399437;
assign t[1256] = 3146;
assign s[1257] = 10396290;
assign t[1257] = 3144;
assign s[1258] = 10393146;
assign t[1258] = 3142;
assign s[1259] = 10390003;
assign t[1259] = 3140;
assign s[1260] = 10386862;
assign t[1260] = 3138;
assign s[1261] = 10383723;
assign t[1261] = 3137;
assign s[1262] = 10380586;
assign t[1262] = 3135;
assign s[1263] = 10377451;
assign t[1263] = 3133;
assign s[1264] = 10374317;
assign t[1264] = 3131;
assign s[1265] = 10371186;
assign t[1265] = 3129;
assign s[1266] = 10368057;
assign t[1266] = 3127;
assign s[1267] = 10364929;
assign t[1267] = 3125;
assign s[1268] = 10361803;
assign t[1268] = 3123;
assign s[1269] = 10358679;
assign t[1269] = 3121;
assign s[1270] = 10355557;
assign t[1270] = 3120;
assign s[1271] = 10352437;
assign t[1271] = 3118;
assign s[1272] = 10349319;
assign t[1272] = 3116;
assign s[1273] = 10346203;
assign t[1273] = 3114;
assign s[1274] = 10343088;
assign t[1274] = 3112;
assign s[1275] = 10339976;
assign t[1275] = 3110;
assign s[1276] = 10336865;
assign t[1276] = 3108;
assign s[1277] = 10333756;
assign t[1277] = 3106;
assign s[1278] = 10330649;
assign t[1278] = 3105;
assign s[1279] = 10327544;
assign t[1279] = 3103;
assign s[1280] = 10324441;
assign t[1280] = 3101;
assign s[1281] = 10321340;
assign t[1281] = 3099;
assign s[1282] = 10318240;
assign t[1282] = 3097;
assign s[1283] = 10315142;
assign t[1283] = 3095;
assign s[1284] = 10312047;
assign t[1284] = 3093;
assign s[1285] = 10308953;
assign t[1285] = 3092;
assign s[1286] = 10305861;
assign t[1286] = 3090;
assign s[1287] = 10302770;
assign t[1287] = 3088;
assign s[1288] = 10299682;
assign t[1288] = 3086;
assign s[1289] = 10296596;
assign t[1289] = 3084;
assign s[1290] = 10293511;
assign t[1290] = 3082;
assign s[1291] = 10290428;
assign t[1291] = 3080;
assign s[1292] = 10287347;
assign t[1292] = 3079;
assign s[1293] = 10284268;
assign t[1293] = 3077;
assign s[1294] = 10281191;
assign t[1294] = 3075;
assign s[1295] = 10278115;
assign t[1295] = 3073;
assign s[1296] = 10275042;
assign t[1296] = 3071;
assign s[1297] = 10271970;
assign t[1297] = 3069;
assign s[1298] = 10268900;
assign t[1298] = 3068;
assign s[1299] = 10265832;
assign t[1299] = 3066;
assign s[1300] = 10262766;
assign t[1300] = 3064;
assign s[1301] = 10259701;
assign t[1301] = 3062;
assign s[1302] = 10256639;
assign t[1302] = 3060;
assign s[1303] = 10253578;
assign t[1303] = 3058;
assign s[1304] = 10250519;
assign t[1304] = 3057;
assign s[1305] = 10247462;
assign t[1305] = 3055;
assign s[1306] = 10244406;
assign t[1306] = 3053;
assign s[1307] = 10241353;
assign t[1307] = 3051;
assign s[1308] = 10238301;
assign t[1308] = 3049;
assign s[1309] = 10235251;
assign t[1309] = 3048;
assign s[1310] = 10232203;
assign t[1310] = 3046;
assign s[1311] = 10229157;
assign t[1311] = 3044;
assign s[1312] = 10226113;
assign t[1312] = 3042;
assign s[1313] = 10223070;
assign t[1313] = 3040;
assign s[1314] = 10220030;
assign t[1314] = 3038;
assign s[1315] = 10216991;
assign t[1315] = 3037;
assign s[1316] = 10213953;
assign t[1316] = 3035;
assign s[1317] = 10210918;
assign t[1317] = 3033;
assign s[1318] = 10207885;
assign t[1318] = 3031;
assign s[1319] = 10204853;
assign t[1319] = 3029;
assign s[1320] = 10201823;
assign t[1320] = 3028;
assign s[1321] = 10198795;
assign t[1321] = 3026;
assign s[1322] = 10195768;
assign t[1322] = 3024;
assign s[1323] = 10192744;
assign t[1323] = 3022;
assign s[1324] = 10189721;
assign t[1324] = 3020;
assign s[1325] = 10186700;
assign t[1325] = 3019;
assign s[1326] = 10183681;
assign t[1326] = 3017;
assign s[1327] = 10180663;
assign t[1327] = 3015;
assign s[1328] = 10177648;
assign t[1328] = 3013;
assign s[1329] = 10174634;
assign t[1329] = 3012;
assign s[1330] = 10171622;
assign t[1330] = 3010;
assign s[1331] = 10168612;
assign t[1331] = 3008;
assign s[1332] = 10165603;
assign t[1332] = 3006;
assign s[1333] = 10162597;
assign t[1333] = 3004;
assign s[1334] = 10159592;
assign t[1334] = 3003;
assign s[1335] = 10156589;
assign t[1335] = 3001;
assign s[1336] = 10153587;
assign t[1336] = 2999;
assign s[1337] = 10150588;
assign t[1337] = 2997;
assign s[1338] = 10147590;
assign t[1338] = 2996;
assign s[1339] = 10144594;
assign t[1339] = 2994;
assign s[1340] = 10141600;
assign t[1340] = 2992;
assign s[1341] = 10138607;
assign t[1341] = 2990;
assign s[1342] = 10135616;
assign t[1342] = 2988;
assign s[1343] = 10132627;
assign t[1343] = 2987;
assign s[1344] = 10129640;
assign t[1344] = 2985;
assign s[1345] = 10126655;
assign t[1345] = 2983;
assign s[1346] = 10123671;
assign t[1346] = 2981;
assign s[1347] = 10120689;
assign t[1347] = 2980;
assign s[1348] = 10117709;
assign t[1348] = 2978;
assign s[1349] = 10114730;
assign t[1349] = 2976;
assign s[1350] = 10111754;
assign t[1350] = 2974;
assign s[1351] = 10108779;
assign t[1351] = 2973;
assign s[1352] = 10105806;
assign t[1352] = 2971;
assign s[1353] = 10102834;
assign t[1353] = 2969;
assign s[1354] = 10099865;
assign t[1354] = 2967;
assign s[1355] = 10096897;
assign t[1355] = 2966;
assign s[1356] = 10093930;
assign t[1356] = 2964;
assign s[1357] = 10090966;
assign t[1357] = 2962;
assign s[1358] = 10088003;
assign t[1358] = 2960;
assign s[1359] = 10085042;
assign t[1359] = 2959;
assign s[1360] = 10082083;
assign t[1360] = 2957;
assign s[1361] = 10079126;
assign t[1361] = 2955;
assign s[1362] = 10076170;
assign t[1362] = 2954;
assign s[1363] = 10073216;
assign t[1363] = 2952;
assign s[1364] = 10070264;
assign t[1364] = 2950;
assign s[1365] = 10067313;
assign t[1365] = 2948;
assign s[1366] = 10064364;
assign t[1366] = 2947;
assign s[1367] = 10061417;
assign t[1367] = 2945;
assign s[1368] = 10058472;
assign t[1368] = 2943;
assign s[1369] = 10055528;
assign t[1369] = 2941;
assign s[1370] = 10052586;
assign t[1370] = 2940;
assign s[1371] = 10049646;
assign t[1371] = 2938;
assign s[1372] = 10046707;
assign t[1372] = 2936;
assign s[1373] = 10043771;
assign t[1373] = 2935;
assign s[1374] = 10040836;
assign t[1374] = 2933;
assign s[1375] = 10037902;
assign t[1375] = 2931;
assign s[1376] = 10034971;
assign t[1376] = 2929;
assign s[1377] = 10032041;
assign t[1377] = 2928;
assign s[1378] = 10029112;
assign t[1378] = 2926;
assign s[1379] = 10026186;
assign t[1379] = 2924;
assign s[1380] = 10023261;
assign t[1380] = 2923;
assign s[1381] = 10020338;
assign t[1381] = 2921;
assign s[1382] = 10017417;
assign t[1382] = 2919;
assign s[1383] = 10014497;
assign t[1383] = 2917;
assign s[1384] = 10011579;
assign t[1384] = 2916;
assign s[1385] = 10008663;
assign t[1385] = 2914;
assign s[1386] = 10005748;
assign t[1386] = 2912;
assign s[1387] = 10002835;
assign t[1387] = 2911;
assign s[1388] = 9999924;
assign t[1388] = 2909;
assign s[1389] = 9997015;
assign t[1389] = 2907;
assign s[1390] = 9994107;
assign t[1390] = 2906;
assign s[1391] = 9991201;
assign t[1391] = 2904;
assign s[1392] = 9988296;
assign t[1392] = 2902;
assign s[1393] = 9985394;
assign t[1393] = 2901;
assign s[1394] = 9982493;
assign t[1394] = 2899;
assign s[1395] = 9979593;
assign t[1395] = 2897;
assign s[1396] = 9976696;
assign t[1396] = 2895;
assign s[1397] = 9973800;
assign t[1397] = 2894;
assign s[1398] = 9970905;
assign t[1398] = 2892;
assign s[1399] = 9968013;
assign t[1399] = 2890;
assign s[1400] = 9965122;
assign t[1400] = 2889;
assign s[1401] = 9962232;
assign t[1401] = 2887;
assign s[1402] = 9959345;
assign t[1402] = 2885;
assign s[1403] = 9956459;
assign t[1403] = 2884;
assign s[1404] = 9953575;
assign t[1404] = 2882;
assign s[1405] = 9950692;
assign t[1405] = 2880;
assign s[1406] = 9947811;
assign t[1406] = 2879;
assign s[1407] = 9944932;
assign t[1407] = 2877;
assign s[1408] = 9942054;
assign t[1408] = 2875;
assign s[1409] = 9939178;
assign t[1409] = 2874;
assign s[1410] = 9936304;
assign t[1410] = 2872;
assign s[1411] = 9933431;
assign t[1411] = 2870;
assign s[1412] = 9930561;
assign t[1412] = 2869;
assign s[1413] = 9927691;
assign t[1413] = 2867;
assign s[1414] = 9924824;
assign t[1414] = 2865;
assign s[1415] = 9921958;
assign t[1415] = 2864;
assign s[1416] = 9919093;
assign t[1416] = 2862;
assign s[1417] = 9916231;
assign t[1417] = 2861;
assign s[1418] = 9913370;
assign t[1418] = 2859;
assign s[1419] = 9910510;
assign t[1419] = 2857;
assign s[1420] = 9907653;
assign t[1420] = 2856;
assign s[1421] = 9904797;
assign t[1421] = 2854;
assign s[1422] = 9901942;
assign t[1422] = 2852;
assign s[1423] = 9899089;
assign t[1423] = 2851;
assign s[1424] = 9896238;
assign t[1424] = 2849;
assign s[1425] = 9893389;
assign t[1425] = 2847;
assign s[1426] = 9890541;
assign t[1426] = 2846;
assign s[1427] = 9887695;
assign t[1427] = 2844;
assign s[1428] = 9884850;
assign t[1428] = 2842;
assign s[1429] = 9882007;
assign t[1429] = 2841;
assign s[1430] = 9879166;
assign t[1430] = 2839;
assign s[1431] = 9876326;
assign t[1431] = 2838;
assign s[1432] = 9873488;
assign t[1432] = 2836;
assign s[1433] = 9870652;
assign t[1433] = 2834;
assign s[1434] = 9867817;
assign t[1434] = 2833;
assign s[1435] = 9864984;
assign t[1435] = 2831;
assign s[1436] = 9862153;
assign t[1436] = 2829;
assign s[1437] = 9859323;
assign t[1437] = 2828;
assign s[1438] = 9856494;
assign t[1438] = 2826;
assign s[1439] = 9853668;
assign t[1439] = 2825;
assign s[1440] = 9850843;
assign t[1440] = 2823;
assign s[1441] = 9848019;
assign t[1441] = 2821;
assign s[1442] = 9845198;
assign t[1442] = 2820;
assign s[1443] = 9842377;
assign t[1443] = 2818;
assign s[1444] = 9839559;
assign t[1444] = 2816;
assign s[1445] = 9836742;
assign t[1445] = 2815;
assign s[1446] = 9833927;
assign t[1446] = 2813;
assign s[1447] = 9831113;
assign t[1447] = 2812;
assign s[1448] = 9828301;
assign t[1448] = 2810;
assign s[1449] = 9825490;
assign t[1449] = 2808;
assign s[1450] = 9822681;
assign t[1450] = 2807;
assign s[1451] = 9819874;
assign t[1451] = 2805;
assign s[1452] = 9817068;
assign t[1452] = 2804;
assign s[1453] = 9814264;
assign t[1453] = 2802;
assign s[1454] = 9811462;
assign t[1454] = 2800;
assign s[1455] = 9808661;
assign t[1455] = 2799;
assign s[1456] = 9805862;
assign t[1456] = 2797;
assign s[1457] = 9803064;
assign t[1457] = 2796;
assign s[1458] = 9800268;
assign t[1458] = 2794;
assign s[1459] = 9797473;
assign t[1459] = 2792;
assign s[1460] = 9794681;
assign t[1460] = 2791;
assign s[1461] = 9791889;
assign t[1461] = 2789;
assign s[1462] = 9789100;
assign t[1462] = 2788;
assign s[1463] = 9786311;
assign t[1463] = 2786;
assign s[1464] = 9783525;
assign t[1464] = 2784;
assign s[1465] = 9780740;
assign t[1465] = 2783;
assign s[1466] = 9777957;
assign t[1466] = 2781;
assign s[1467] = 9775175;
assign t[1467] = 2780;
assign s[1468] = 9772395;
assign t[1468] = 2778;
assign s[1469] = 9769616;
assign t[1469] = 2777;
assign s[1470] = 9766839;
assign t[1470] = 2775;
assign s[1471] = 9764063;
assign t[1471] = 2773;
assign s[1472] = 9761290;
assign t[1472] = 2772;
assign s[1473] = 9758517;
assign t[1473] = 2770;
assign s[1474] = 9755747;
assign t[1474] = 2769;
assign s[1475] = 9752977;
assign t[1475] = 2767;
assign s[1476] = 9750210;
assign t[1476] = 2766;
assign s[1477] = 9747444;
assign t[1477] = 2764;
assign s[1478] = 9744679;
assign t[1478] = 2762;
assign s[1479] = 9741916;
assign t[1479] = 2761;
assign s[1480] = 9739155;
assign t[1480] = 2759;
assign s[1481] = 9736395;
assign t[1481] = 2758;
assign s[1482] = 9733637;
assign t[1482] = 2756;
assign s[1483] = 9730881;
assign t[1483] = 2755;
assign s[1484] = 9728126;
assign t[1484] = 2753;
assign s[1485] = 9725372;
assign t[1485] = 2751;
assign s[1486] = 9722620;
assign t[1486] = 2750;
assign s[1487] = 9719870;
assign t[1487] = 2748;
assign s[1488] = 9717121;
assign t[1488] = 2747;
assign s[1489] = 9714374;
assign t[1489] = 2745;
assign s[1490] = 9711628;
assign t[1490] = 2744;
assign s[1491] = 9708884;
assign t[1491] = 2742;
assign s[1492] = 9706141;
assign t[1492] = 2741;
assign s[1493] = 9703400;
assign t[1493] = 2739;
assign s[1494] = 9700660;
assign t[1494] = 2737;
assign s[1495] = 9697923;
assign t[1495] = 2736;
assign s[1496] = 9695186;
assign t[1496] = 2734;
assign s[1497] = 9692451;
assign t[1497] = 2733;
assign s[1498] = 9689718;
assign t[1498] = 2731;
assign s[1499] = 9686986;
assign t[1499] = 2730;
assign s[1500] = 9684256;
assign t[1500] = 2728;
assign s[1501] = 9681527;
assign t[1501] = 2727;
assign s[1502] = 9678800;
assign t[1502] = 2725;
assign s[1503] = 9676074;
assign t[1503] = 2724;
assign s[1504] = 9673350;
assign t[1504] = 2722;
assign s[1505] = 9670627;
assign t[1505] = 2721;
assign s[1506] = 9667906;
assign t[1506] = 2719;
assign s[1507] = 9665187;
assign t[1507] = 2717;
assign s[1508] = 9662469;
assign t[1508] = 2716;
assign s[1509] = 9659752;
assign t[1509] = 2714;
assign s[1510] = 9657038;
assign t[1510] = 2713;
assign s[1511] = 9654324;
assign t[1511] = 2711;
assign s[1512] = 9651612;
assign t[1512] = 2710;
assign s[1513] = 9648902;
assign t[1513] = 2708;
assign s[1514] = 9646193;
assign t[1514] = 2707;
assign s[1515] = 9643486;
assign t[1515] = 2705;
assign s[1516] = 9640780;
assign t[1516] = 2704;
assign s[1517] = 9638076;
assign t[1517] = 2702;
assign s[1518] = 9635373;
assign t[1518] = 2701;
assign s[1519] = 9632672;
assign t[1519] = 2699;
assign s[1520] = 9629972;
assign t[1520] = 2698;
assign s[1521] = 9627274;
assign t[1521] = 2696;
assign s[1522] = 9624577;
assign t[1522] = 2695;
assign s[1523] = 9621882;
assign t[1523] = 2693;
assign s[1524] = 9619188;
assign t[1524] = 2692;
assign s[1525] = 9616496;
assign t[1525] = 2690;
assign s[1526] = 9613805;
assign t[1526] = 2689;
assign s[1527] = 9611116;
assign t[1527] = 2687;
assign s[1528] = 9608428;
assign t[1528] = 2686;
assign s[1529] = 9605742;
assign t[1529] = 2684;
assign s[1530] = 9603057;
assign t[1530] = 2683;
assign s[1531] = 9600374;
assign t[1531] = 2681;
assign s[1532] = 9597693;
assign t[1532] = 2680;
assign s[1533] = 9595012;
assign t[1533] = 2678;
assign s[1534] = 9592334;
assign t[1534] = 2677;
assign s[1535] = 9589657;
assign t[1535] = 2675;
assign s[1536] = 9586981;
assign t[1536] = 2674;
assign s[1537] = 9584307;
assign t[1537] = 2672;
assign s[1538] = 9581634;
assign t[1538] = 2671;
assign s[1539] = 9578963;
assign t[1539] = 2669;
assign s[1540] = 9576293;
assign t[1540] = 2668;
assign s[1541] = 9573625;
assign t[1541] = 2666;
assign s[1542] = 9570958;
assign t[1542] = 2665;
assign s[1543] = 9568293;
assign t[1543] = 2663;
assign s[1544] = 9565629;
assign t[1544] = 2662;
assign s[1545] = 9562967;
assign t[1545] = 2660;
assign s[1546] = 9560306;
assign t[1546] = 2659;
assign s[1547] = 9557647;
assign t[1547] = 2657;
assign s[1548] = 9554989;
assign t[1548] = 2656;
assign s[1549] = 9552332;
assign t[1549] = 2654;
assign s[1550] = 9549677;
assign t[1550] = 2653;
assign s[1551] = 9547024;
assign t[1551] = 2651;
assign s[1552] = 9544372;
assign t[1552] = 2650;
assign s[1553] = 9541722;
assign t[1553] = 2649;
assign s[1554] = 9539073;
assign t[1554] = 2647;
assign s[1555] = 9536425;
assign t[1555] = 2646;
assign s[1556] = 9533779;
assign t[1556] = 2644;
assign s[1557] = 9531134;
assign t[1557] = 2643;
assign s[1558] = 9528491;
assign t[1558] = 2641;
assign s[1559] = 9525850;
assign t[1559] = 2640;
assign s[1560] = 9523209;
assign t[1560] = 2638;
assign s[1561] = 9520571;
assign t[1561] = 2637;
assign s[1562] = 9517933;
assign t[1562] = 2635;
assign s[1563] = 9515298;
assign t[1563] = 2634;
assign s[1564] = 9512663;
assign t[1564] = 2632;
assign s[1565] = 9510030;
assign t[1565] = 2631;
assign s[1566] = 9507399;
assign t[1566] = 2629;
assign s[1567] = 9504769;
assign t[1567] = 2628;
assign s[1568] = 9502140;
assign t[1568] = 2627;
assign s[1569] = 9499513;
assign t[1569] = 2625;
assign s[1570] = 9496888;
assign t[1570] = 2624;
assign s[1571] = 9494263;
assign t[1571] = 2622;
assign s[1572] = 9491641;
assign t[1572] = 2621;
assign s[1573] = 9489019;
assign t[1573] = 2619;
assign s[1574] = 9486400;
assign t[1574] = 2618;
assign s[1575] = 9483781;
assign t[1575] = 2616;
assign s[1576] = 9481164;
assign t[1576] = 2615;
assign s[1577] = 9478549;
assign t[1577] = 2614;
assign s[1578] = 9475935;
assign t[1578] = 2612;
assign s[1579] = 9473322;
assign t[1579] = 2611;
assign s[1580] = 9470711;
assign t[1580] = 2609;
assign s[1581] = 9468101;
assign t[1581] = 2608;
assign s[1582] = 9465493;
assign t[1582] = 2606;
assign s[1583] = 9462886;
assign t[1583] = 2605;
assign s[1584] = 9460281;
assign t[1584] = 2603;
assign s[1585] = 9457677;
assign t[1585] = 2602;
assign s[1586] = 9455074;
assign t[1586] = 2601;
assign s[1587] = 9452473;
assign t[1587] = 2599;
assign s[1588] = 9449873;
assign t[1588] = 2598;
assign s[1589] = 9447275;
assign t[1589] = 2596;
assign s[1590] = 9444678;
assign t[1590] = 2595;
assign s[1591] = 9442083;
assign t[1591] = 2593;
assign s[1592] = 9439489;
assign t[1592] = 2592;
assign s[1593] = 9436896;
assign t[1593] = 2591;
assign s[1594] = 9434305;
assign t[1594] = 2589;
assign s[1595] = 9431715;
assign t[1595] = 2588;
assign s[1596] = 9429127;
assign t[1596] = 2586;
assign s[1597] = 9426540;
assign t[1597] = 2585;
assign s[1598] = 9423955;
assign t[1598] = 2584;
assign s[1599] = 9421371;
assign t[1599] = 2582;
assign s[1600] = 9418788;
assign t[1600] = 2581;
assign s[1601] = 9416207;
assign t[1601] = 2579;
assign s[1602] = 9413627;
assign t[1602] = 2578;
assign s[1603] = 9411049;
assign t[1603] = 2576;
assign s[1604] = 9408472;
assign t[1604] = 2575;
assign s[1605] = 9405896;
assign t[1605] = 2574;
assign s[1606] = 9403322;
assign t[1606] = 2572;
assign s[1607] = 9400750;
assign t[1607] = 2571;
assign s[1608] = 9398178;
assign t[1608] = 2569;
assign s[1609] = 9395608;
assign t[1609] = 2568;
assign s[1610] = 9393040;
assign t[1610] = 2567;
assign s[1611] = 9390473;
assign t[1611] = 2565;
assign s[1612] = 9387907;
assign t[1612] = 2564;
assign s[1613] = 9385343;
assign t[1613] = 2562;
assign s[1614] = 9382780;
assign t[1614] = 2561;
assign s[1615] = 9380218;
assign t[1615] = 2560;
assign s[1616] = 9377658;
assign t[1616] = 2558;
assign s[1617] = 9375099;
assign t[1617] = 2557;
assign s[1618] = 9372542;
assign t[1618] = 2555;
assign s[1619] = 9369986;
assign t[1619] = 2554;
assign s[1620] = 9367432;
assign t[1620] = 2553;
assign s[1621] = 9364879;
assign t[1621] = 2551;
assign s[1622] = 9362327;
assign t[1622] = 2550;
assign s[1623] = 9359777;
assign t[1623] = 2548;
assign s[1624] = 9357228;
assign t[1624] = 2547;
assign s[1625] = 9354680;
assign t[1625] = 2546;
assign s[1626] = 9352134;
assign t[1626] = 2544;
assign s[1627] = 9349589;
assign t[1627] = 2543;
assign s[1628] = 9347046;
assign t[1628] = 2542;
assign s[1629] = 9344504;
assign t[1629] = 2540;
assign s[1630] = 9341963;
assign t[1630] = 2539;
assign s[1631] = 9339424;
assign t[1631] = 2537;
assign s[1632] = 9336886;
assign t[1632] = 2536;
assign s[1633] = 9334349;
assign t[1633] = 2535;
assign s[1634] = 9331814;
assign t[1634] = 2533;
assign s[1635] = 9329280;
assign t[1635] = 2532;
assign s[1636] = 9326748;
assign t[1636] = 2531;
assign s[1637] = 9324217;
assign t[1637] = 2529;
assign s[1638] = 9321687;
assign t[1638] = 2528;
assign s[1639] = 9319159;
assign t[1639] = 2526;
assign s[1640] = 9316632;
assign t[1640] = 2525;
assign s[1641] = 9314107;
assign t[1641] = 2524;
assign s[1642] = 9311583;
assign t[1642] = 2522;
assign s[1643] = 9309060;
assign t[1643] = 2521;
assign s[1644] = 9306538;
assign t[1644] = 2520;
assign s[1645] = 9304018;
assign t[1645] = 2518;
assign s[1646] = 9301500;
assign t[1646] = 2517;
assign s[1647] = 9298982;
assign t[1647] = 2515;
assign s[1648] = 9296466;
assign t[1648] = 2514;
assign s[1649] = 9293952;
assign t[1649] = 2513;
assign s[1650] = 9291439;
assign t[1650] = 2511;
assign s[1651] = 9288927;
assign t[1651] = 2510;
assign s[1652] = 9286416;
assign t[1652] = 2509;
assign s[1653] = 9283907;
assign t[1653] = 2507;
assign s[1654] = 9281399;
assign t[1654] = 2506;
assign s[1655] = 9278893;
assign t[1655] = 2505;
assign s[1656] = 9276388;
assign t[1656] = 2503;
assign s[1657] = 9273884;
assign t[1657] = 2502;
assign s[1658] = 9271381;
assign t[1658] = 2501;
assign s[1659] = 9268880;
assign t[1659] = 2499;
assign s[1660] = 9266381;
assign t[1660] = 2498;
assign s[1661] = 9263882;
assign t[1661] = 2497;
assign s[1662] = 9261385;
assign t[1662] = 2495;
assign s[1663] = 9258890;
assign t[1663] = 2494;
assign s[1664] = 9256395;
assign t[1664] = 2492;
assign s[1665] = 9253902;
assign t[1665] = 2491;
assign s[1666] = 9251411;
assign t[1666] = 2490;
assign s[1667] = 9248920;
assign t[1667] = 2488;
assign s[1668] = 9246432;
assign t[1668] = 2487;
assign s[1669] = 9243944;
assign t[1669] = 2486;
assign s[1670] = 9241458;
assign t[1670] = 2484;
assign s[1671] = 9238973;
assign t[1671] = 2483;
assign s[1672] = 9236489;
assign t[1672] = 2482;
assign s[1673] = 9234007;
assign t[1673] = 2480;
assign s[1674] = 9231526;
assign t[1674] = 2479;
assign s[1675] = 9229046;
assign t[1675] = 2478;
assign s[1676] = 9226568;
assign t[1676] = 2476;
assign s[1677] = 9224091;
assign t[1677] = 2475;
assign s[1678] = 9221616;
assign t[1678] = 2474;
assign s[1679] = 9219141;
assign t[1679] = 2472;
assign s[1680] = 9216668;
assign t[1680] = 2471;
assign s[1681] = 9214197;
assign t[1681] = 2470;
assign s[1682] = 9211726;
assign t[1682] = 2468;
assign s[1683] = 9209257;
assign t[1683] = 2467;
assign s[1684] = 9206790;
assign t[1684] = 2466;
assign s[1685] = 9204323;
assign t[1685] = 2465;
assign s[1686] = 9201858;
assign t[1686] = 2463;
assign s[1687] = 9199395;
assign t[1687] = 2462;
assign s[1688] = 9196932;
assign t[1688] = 2461;
assign s[1689] = 9194471;
assign t[1689] = 2459;
assign s[1690] = 9192012;
assign t[1690] = 2458;
assign s[1691] = 9189553;
assign t[1691] = 2457;
assign s[1692] = 9187096;
assign t[1692] = 2455;
assign s[1693] = 9184640;
assign t[1693] = 2454;
assign s[1694] = 9182186;
assign t[1694] = 2453;
assign s[1695] = 9179733;
assign t[1695] = 2451;
assign s[1696] = 9177281;
assign t[1696] = 2450;
assign s[1697] = 9174830;
assign t[1697] = 2449;
assign s[1698] = 9172381;
assign t[1698] = 2447;
assign s[1699] = 9169933;
assign t[1699] = 2446;
assign s[1700] = 9167487;
assign t[1700] = 2445;
assign s[1701] = 9165041;
assign t[1701] = 2444;
assign s[1702] = 9162597;
assign t[1702] = 2442;
assign s[1703] = 9160155;
assign t[1703] = 2441;
assign s[1704] = 9157713;
assign t[1704] = 2440;
assign s[1705] = 9155273;
assign t[1705] = 2438;
assign s[1706] = 9152834;
assign t[1706] = 2437;
assign s[1707] = 9150397;
assign t[1707] = 2436;
assign s[1708] = 9147960;
assign t[1708] = 2434;
assign s[1709] = 9145526;
assign t[1709] = 2433;
assign s[1710] = 9143092;
assign t[1710] = 2432;
assign s[1711] = 9140660;
assign t[1711] = 2431;
assign s[1712] = 9138229;
assign t[1712] = 2429;
assign s[1713] = 9135799;
assign t[1713] = 2428;
assign s[1714] = 9133370;
assign t[1714] = 2427;
assign s[1715] = 9130943;
assign t[1715] = 2425;
assign s[1716] = 9128517;
assign t[1716] = 2424;
assign s[1717] = 9126093;
assign t[1717] = 2423;
assign s[1718] = 9123670;
assign t[1718] = 2421;
assign s[1719] = 9121248;
assign t[1719] = 2420;
assign s[1720] = 9118827;
assign t[1720] = 2419;
assign s[1721] = 9116407;
assign t[1721] = 2418;
assign s[1722] = 9113989;
assign t[1722] = 2416;
assign s[1723] = 9111572;
assign t[1723] = 2415;
assign s[1724] = 9109157;
assign t[1724] = 2414;
assign s[1725] = 9106743;
assign t[1725] = 2413;
assign s[1726] = 9104330;
assign t[1726] = 2411;
assign s[1727] = 9101918;
assign t[1727] = 2410;
assign s[1728] = 9099507;
assign t[1728] = 2409;
assign s[1729] = 9097098;
assign t[1729] = 2407;
assign s[1730] = 9094690;
assign t[1730] = 2406;
assign s[1731] = 9092284;
assign t[1731] = 2405;
assign s[1732] = 9089878;
assign t[1732] = 2404;
assign s[1733] = 9087474;
assign t[1733] = 2402;
assign s[1734] = 9085071;
assign t[1734] = 2401;
assign s[1735] = 9082670;
assign t[1735] = 2400;
assign s[1736] = 9080269;
assign t[1736] = 2399;
assign s[1737] = 9077870;
assign t[1737] = 2397;
assign s[1738] = 9075473;
assign t[1738] = 2396;
assign s[1739] = 9073076;
assign t[1739] = 2395;
assign s[1740] = 9070681;
assign t[1740] = 2393;
assign s[1741] = 9068287;
assign t[1741] = 2392;
assign s[1742] = 9065894;
assign t[1742] = 2391;
assign s[1743] = 9063503;
assign t[1743] = 2390;
assign s[1744] = 9061113;
assign t[1744] = 2388;
assign s[1745] = 9058724;
assign t[1745] = 2387;
assign s[1746] = 9056336;
assign t[1746] = 2386;
assign s[1747] = 9053950;
assign t[1747] = 2385;
assign s[1748] = 9051565;
assign t[1748] = 2383;
assign s[1749] = 9049181;
assign t[1749] = 2382;
assign s[1750] = 9046798;
assign t[1750] = 2381;
assign s[1751] = 9044417;
assign t[1751] = 2380;
assign s[1752] = 9042037;
assign t[1752] = 2378;
assign s[1753] = 9039658;
assign t[1753] = 2377;
assign s[1754] = 9037280;
assign t[1754] = 2376;
assign s[1755] = 9034904;
assign t[1755] = 2375;
assign s[1756] = 9032529;
assign t[1756] = 2373;
assign s[1757] = 9030155;
assign t[1757] = 2372;
assign s[1758] = 9027782;
assign t[1758] = 2371;
assign s[1759] = 9025411;
assign t[1759] = 2370;
assign s[1760] = 9023041;
assign t[1760] = 2368;
assign s[1761] = 9020672;
assign t[1761] = 2367;
assign s[1762] = 9018304;
assign t[1762] = 2366;
assign s[1763] = 9015938;
assign t[1763] = 2365;
assign s[1764] = 9013573;
assign t[1764] = 2363;
assign s[1765] = 9011209;
assign t[1765] = 2362;
assign s[1766] = 9008846;
assign t[1766] = 2361;
assign s[1767] = 9006485;
assign t[1767] = 2360;
assign s[1768] = 9004125;
assign t[1768] = 2358;
assign s[1769] = 9001766;
assign t[1769] = 2357;
assign s[1770] = 8999408;
assign t[1770] = 2356;
assign s[1771] = 8997052;
assign t[1771] = 2355;
assign s[1772] = 8994696;
assign t[1772] = 2354;
assign s[1773] = 8992342;
assign t[1773] = 2352;
assign s[1774] = 8989989;
assign t[1774] = 2351;
assign s[1775] = 8987638;
assign t[1775] = 2350;
assign s[1776] = 8985288;
assign t[1776] = 2349;
assign s[1777] = 8982938;
assign t[1777] = 2347;
assign s[1778] = 8980591;
assign t[1778] = 2346;
assign s[1779] = 8978244;
assign t[1779] = 2345;
assign s[1780] = 8975899;
assign t[1780] = 2344;
assign s[1781] = 8973554;
assign t[1781] = 2342;
assign s[1782] = 8971211;
assign t[1782] = 2341;
assign s[1783] = 8968870;
assign t[1783] = 2340;
assign s[1784] = 8966529;
assign t[1784] = 2339;
assign s[1785] = 8964190;
assign t[1785] = 2338;
assign s[1786] = 8961852;
assign t[1786] = 2336;
assign s[1787] = 8959515;
assign t[1787] = 2335;
assign s[1788] = 8957179;
assign t[1788] = 2334;
assign s[1789] = 8954845;
assign t[1789] = 2333;
assign s[1790] = 8952512;
assign t[1790] = 2331;
assign s[1791] = 8950180;
assign t[1791] = 2330;
assign s[1792] = 8947849;
assign t[1792] = 2329;
assign s[1793] = 8945519;
assign t[1793] = 2328;
assign s[1794] = 8943191;
assign t[1794] = 2327;
assign s[1795] = 8940864;
assign t[1795] = 2325;
assign s[1796] = 8938538;
assign t[1796] = 2324;
assign s[1797] = 8936213;
assign t[1797] = 2323;
assign s[1798] = 8933890;
assign t[1798] = 2322;
assign s[1799] = 8931567;
assign t[1799] = 2321;
assign s[1800] = 8929246;
assign t[1800] = 2319;
assign s[1801] = 8926926;
assign t[1801] = 2318;
assign s[1802] = 8924608;
assign t[1802] = 2317;
assign s[1803] = 8922290;
assign t[1803] = 2316;
assign s[1804] = 8919974;
assign t[1804] = 2315;
assign s[1805] = 8917659;
assign t[1805] = 2313;
assign s[1806] = 8915345;
assign t[1806] = 2312;
assign s[1807] = 8913032;
assign t[1807] = 2311;
assign s[1808] = 8910721;
assign t[1808] = 2310;
assign s[1809] = 8908411;
assign t[1809] = 2309;
assign s[1810] = 8906102;
assign t[1810] = 2307;
assign s[1811] = 8903794;
assign t[1811] = 2306;
assign s[1812] = 8901487;
assign t[1812] = 2305;
assign s[1813] = 8899181;
assign t[1813] = 2304;
assign s[1814] = 8896877;
assign t[1814] = 2303;
assign s[1815] = 8894574;
assign t[1815] = 2301;
assign s[1816] = 8892272;
assign t[1816] = 2300;
assign s[1817] = 8889971;
assign t[1817] = 2299;
assign s[1818] = 8887672;
assign t[1818] = 2298;
assign s[1819] = 8885374;
assign t[1819] = 2297;
assign s[1820] = 8883076;
assign t[1820] = 2295;
assign s[1821] = 8880780;
assign t[1821] = 2294;
assign s[1822] = 8878486;
assign t[1822] = 2293;
assign s[1823] = 8876192;
assign t[1823] = 2292;
assign s[1824] = 8873900;
assign t[1824] = 2291;
assign s[1825] = 8871609;
assign t[1825] = 2290;
assign s[1826] = 8869318;
assign t[1826] = 2288;
assign s[1827] = 8867030;
assign t[1827] = 2287;
assign s[1828] = 8864742;
assign t[1828] = 2286;
assign s[1829] = 8862455;
assign t[1829] = 2285;
assign s[1830] = 8860170;
assign t[1830] = 2284;
assign s[1831] = 8857886;
assign t[1831] = 2282;
assign s[1832] = 8855603;
assign t[1832] = 2281;
assign s[1833] = 8853321;
assign t[1833] = 2280;
assign s[1834] = 8851041;
assign t[1834] = 2279;
assign s[1835] = 8848761;
assign t[1835] = 2278;
assign s[1836] = 8846483;
assign t[1836] = 2277;
assign s[1837] = 8844206;
assign t[1837] = 2275;
assign s[1838] = 8841930;
assign t[1838] = 2274;
assign s[1839] = 8839655;
assign t[1839] = 2273;
assign s[1840] = 8837382;
assign t[1840] = 2272;
assign s[1841] = 8835109;
assign t[1841] = 2271;
assign s[1842] = 8832838;
assign t[1842] = 2270;
assign s[1843] = 8830568;
assign t[1843] = 2268;
assign s[1844] = 8828299;
assign t[1844] = 2267;
assign s[1845] = 8826031;
assign t[1845] = 2266;
assign s[1846] = 8823765;
assign t[1846] = 2265;
assign s[1847] = 8821499;
assign t[1847] = 2264;
assign s[1848] = 8819235;
assign t[1848] = 2263;
assign s[1849] = 8816972;
assign t[1849] = 2261;
assign s[1850] = 8814710;
assign t[1850] = 2260;
assign s[1851] = 8812449;
assign t[1851] = 2259;
assign s[1852] = 8810190;
assign t[1852] = 2258;
assign s[1853] = 8807931;
assign t[1853] = 2257;
assign s[1854] = 8805674;
assign t[1854] = 2256;
assign s[1855] = 8803418;
assign t[1855] = 2254;
assign s[1856] = 8801163;
assign t[1856] = 2253;
assign s[1857] = 8798909;
assign t[1857] = 2252;
assign s[1858] = 8796656;
assign t[1858] = 2251;
assign s[1859] = 8794405;
assign t[1859] = 2250;
assign s[1860] = 8792154;
assign t[1860] = 2249;
assign s[1861] = 8789905;
assign t[1861] = 2248;
assign s[1862] = 8787657;
assign t[1862] = 2246;
assign s[1863] = 8785410;
assign t[1863] = 2245;
assign s[1864] = 8783165;
assign t[1864] = 2244;
assign s[1865] = 8780920;
assign t[1865] = 2243;
assign s[1866] = 8778676;
assign t[1866] = 2242;
assign s[1867] = 8776434;
assign t[1867] = 2241;
assign s[1868] = 8774193;
assign t[1868] = 2240;
assign s[1869] = 8771953;
assign t[1869] = 2238;
assign s[1870] = 8769714;
assign t[1870] = 2237;
assign s[1871] = 8767476;
assign t[1871] = 2236;
assign s[1872] = 8765240;
assign t[1872] = 2235;
assign s[1873] = 8763004;
assign t[1873] = 2234;
assign s[1874] = 8760770;
assign t[1874] = 2233;
assign s[1875] = 8758537;
assign t[1875] = 2232;
assign s[1876] = 8756305;
assign t[1876] = 2230;
assign s[1877] = 8754074;
assign t[1877] = 2229;
assign s[1878] = 8751844;
assign t[1878] = 2228;
assign s[1879] = 8749615;
assign t[1879] = 2227;
assign s[1880] = 8747388;
assign t[1880] = 2226;
assign s[1881] = 8745162;
assign t[1881] = 2225;
assign s[1882] = 8742936;
assign t[1882] = 2224;
assign s[1883] = 8740712;
assign t[1883] = 2222;
assign s[1884] = 8738489;
assign t[1884] = 2221;
assign s[1885] = 8736267;
assign t[1885] = 2220;
assign s[1886] = 8734047;
assign t[1886] = 2219;
assign s[1887] = 8731827;
assign t[1887] = 2218;
assign s[1888] = 8729609;
assign t[1888] = 2217;
assign s[1889] = 8727391;
assign t[1889] = 2216;
assign s[1890] = 8725175;
assign t[1890] = 2215;
assign s[1891] = 8722960;
assign t[1891] = 2213;
assign s[1892] = 8720746;
assign t[1892] = 2212;
assign s[1893] = 8718533;
assign t[1893] = 2211;
assign s[1894] = 8716322;
assign t[1894] = 2210;
assign s[1895] = 8714111;
assign t[1895] = 2209;
assign s[1896] = 8711902;
assign t[1896] = 2208;
assign s[1897] = 8709693;
assign t[1897] = 2207;
assign s[1898] = 8707486;
assign t[1898] = 2206;
assign s[1899] = 8705280;
assign t[1899] = 2204;
assign s[1900] = 8703075;
assign t[1900] = 2203;
assign s[1901] = 8700871;
assign t[1901] = 2202;
assign s[1902] = 8698668;
assign t[1902] = 2201;
assign s[1903] = 8696467;
assign t[1903] = 2200;
assign s[1904] = 8694266;
assign t[1904] = 2199;
assign s[1905] = 8692067;
assign t[1905] = 2198;
assign s[1906] = 8689868;
assign t[1906] = 2197;
assign s[1907] = 8687671;
assign t[1907] = 2196;
assign s[1908] = 8685475;
assign t[1908] = 2194;
assign s[1909] = 8683280;
assign t[1909] = 2193;
assign s[1910] = 8681086;
assign t[1910] = 2192;
assign s[1911] = 8678894;
assign t[1911] = 2191;
assign s[1912] = 8676702;
assign t[1912] = 2190;
assign s[1913] = 8674511;
assign t[1913] = 2189;
assign s[1914] = 8672322;
assign t[1914] = 2188;
assign s[1915] = 8670134;
assign t[1915] = 2187;
assign s[1916] = 8667946;
assign t[1916] = 2186;
assign s[1917] = 8665760;
assign t[1917] = 2185;
assign s[1918] = 8663575;
assign t[1918] = 2183;
assign s[1919] = 8661391;
assign t[1919] = 2182;
assign s[1920] = 8659209;
assign t[1920] = 2181;
assign s[1921] = 8657027;
assign t[1921] = 2180;
assign s[1922] = 8654846;
assign t[1922] = 2179;
assign s[1923] = 8652667;
assign t[1923] = 2178;
assign s[1924] = 8650488;
assign t[1924] = 2177;
assign s[1925] = 8648311;
assign t[1925] = 2176;
assign s[1926] = 8646135;
assign t[1926] = 2175;
assign s[1927] = 8643960;
assign t[1927] = 2174;
assign s[1928] = 8641786;
assign t[1928] = 2172;
assign s[1929] = 8639613;
assign t[1929] = 2171;
assign s[1930] = 8637441;
assign t[1930] = 2170;
assign s[1931] = 8635270;
assign t[1931] = 2169;
assign s[1932] = 8633100;
assign t[1932] = 2168;
assign s[1933] = 8630932;
assign t[1933] = 2167;
assign s[1934] = 8628764;
assign t[1934] = 2166;
assign s[1935] = 8626598;
assign t[1935] = 2165;
assign s[1936] = 8624433;
assign t[1936] = 2164;
assign s[1937] = 8622268;
assign t[1937] = 2163;
assign s[1938] = 8620105;
assign t[1938] = 2162;
assign s[1939] = 8617943;
assign t[1939] = 2160;
assign s[1940] = 8615782;
assign t[1940] = 2159;
assign s[1941] = 8613622;
assign t[1941] = 2158;
assign s[1942] = 8611464;
assign t[1942] = 2157;
assign s[1943] = 8609306;
assign t[1943] = 2156;
assign s[1944] = 8607149;
assign t[1944] = 2155;
assign s[1945] = 8604994;
assign t[1945] = 2154;
assign s[1946] = 8602839;
assign t[1946] = 2153;
assign s[1947] = 8600686;
assign t[1947] = 2152;
assign s[1948] = 8598533;
assign t[1948] = 2151;
assign s[1949] = 8596382;
assign t[1949] = 2150;
assign s[1950] = 8594232;
assign t[1950] = 2149;
assign s[1951] = 8592083;
assign t[1951] = 2148;
assign s[1952] = 8589935;
assign t[1952] = 2146;
assign s[1953] = 8587788;
assign t[1953] = 2145;
assign s[1954] = 8585642;
assign t[1954] = 2144;
assign s[1955] = 8583497;
assign t[1955] = 2143;
assign s[1956] = 8581354;
assign t[1956] = 2142;
assign s[1957] = 8579211;
assign t[1957] = 2141;
assign s[1958] = 8577069;
assign t[1958] = 2140;
assign s[1959] = 8574929;
assign t[1959] = 2139;
assign s[1960] = 8572789;
assign t[1960] = 2138;
assign s[1961] = 8570651;
assign t[1961] = 2137;
assign s[1962] = 8568514;
assign t[1962] = 2136;
assign s[1963] = 8566377;
assign t[1963] = 2135;
assign s[1964] = 8564242;
assign t[1964] = 2134;
assign s[1965] = 8562108;
assign t[1965] = 2133;
assign s[1966] = 8559975;
assign t[1966] = 2131;
assign s[1967] = 8557843;
assign t[1967] = 2130;
assign s[1968] = 8555712;
assign t[1968] = 2129;
assign s[1969] = 8553582;
assign t[1969] = 2128;
assign s[1970] = 8551453;
assign t[1970] = 2127;
assign s[1971] = 8549326;
assign t[1971] = 2126;
assign s[1972] = 8547199;
assign t[1972] = 2125;
assign s[1973] = 8545073;
assign t[1973] = 2124;
assign s[1974] = 8542949;
assign t[1974] = 2123;
assign s[1975] = 8540825;
assign t[1975] = 2122;
assign s[1976] = 8538703;
assign t[1976] = 2121;
assign s[1977] = 8536581;
assign t[1977] = 2120;
assign s[1978] = 8534461;
assign t[1978] = 2119;
assign s[1979] = 8532342;
assign t[1979] = 2118;
assign s[1980] = 8530223;
assign t[1980] = 2117;
assign s[1981] = 8528106;
assign t[1981] = 2116;
assign s[1982] = 8525990;
assign t[1982] = 2115;
assign s[1983] = 8523875;
assign t[1983] = 2114;
assign s[1984] = 8521761;
assign t[1984] = 2113;
assign s[1985] = 8519648;
assign t[1985] = 2111;
assign s[1986] = 8517536;
assign t[1986] = 2110;
assign s[1987] = 8515425;
assign t[1987] = 2109;
assign s[1988] = 8513315;
assign t[1988] = 2108;
assign s[1989] = 8511206;
assign t[1989] = 2107;
assign s[1990] = 8509099;
assign t[1990] = 2106;
assign s[1991] = 8506992;
assign t[1991] = 2105;
assign s[1992] = 8504886;
assign t[1992] = 2104;
assign s[1993] = 8502781;
assign t[1993] = 2103;
assign s[1994] = 8500678;
assign t[1994] = 2102;
assign s[1995] = 8498575;
assign t[1995] = 2101;
assign s[1996] = 8496474;
assign t[1996] = 2100;
assign s[1997] = 8494373;
assign t[1997] = 2099;
assign s[1998] = 8492274;
assign t[1998] = 2098;
assign s[1999] = 8490175;
assign t[1999] = 2097;
assign s[2000] = 8488078;
assign t[2000] = 2096;
assign s[2001] = 8485982;
assign t[2001] = 2095;
assign s[2002] = 8483886;
assign t[2002] = 2094;
assign s[2003] = 8481792;
assign t[2003] = 2093;
assign s[2004] = 8479699;
assign t[2004] = 2092;
assign s[2005] = 8477607;
assign t[2005] = 2091;
assign s[2006] = 8475516;
assign t[2006] = 2090;
assign s[2007] = 8473425;
assign t[2007] = 2089;
assign s[2008] = 8471336;
assign t[2008] = 2088;
assign s[2009] = 8469248;
assign t[2009] = 2087;
assign s[2010] = 8467161;
assign t[2010] = 2086;
assign s[2011] = 8465075;
assign t[2011] = 2084;
assign s[2012] = 8462990;
assign t[2012] = 2083;
assign s[2013] = 8460906;
assign t[2013] = 2082;
assign s[2014] = 8458823;
assign t[2014] = 2081;
assign s[2015] = 8456741;
assign t[2015] = 2080;
assign s[2016] = 8454660;
assign t[2016] = 2079;
assign s[2017] = 8452581;
assign t[2017] = 2078;
assign s[2018] = 8450502;
assign t[2018] = 2077;
assign s[2019] = 8448424;
assign t[2019] = 2076;
assign s[2020] = 8446347;
assign t[2020] = 2075;
assign s[2021] = 8444271;
assign t[2021] = 2074;
assign s[2022] = 8442197;
assign t[2022] = 2073;
assign s[2023] = 8440123;
assign t[2023] = 2072;
assign s[2024] = 8438050;
assign t[2024] = 2071;
assign s[2025] = 8435978;
assign t[2025] = 2070;
assign s[2026] = 8433908;
assign t[2026] = 2069;
assign s[2027] = 8431838;
assign t[2027] = 2068;
assign s[2028] = 8429769;
assign t[2028] = 2067;
assign s[2029] = 8427702;
assign t[2029] = 2066;
assign s[2030] = 8425635;
assign t[2030] = 2065;
assign s[2031] = 8423569;
assign t[2031] = 2064;
assign s[2032] = 8421505;
assign t[2032] = 2063;
assign s[2033] = 8419441;
assign t[2033] = 2062;
assign s[2034] = 8417379;
assign t[2034] = 2061;
assign s[2035] = 8415317;
assign t[2035] = 2060;
assign s[2036] = 8413257;
assign t[2036] = 2059;
assign s[2037] = 8411197;
assign t[2037] = 2058;
assign s[2038] = 8409138;
assign t[2038] = 2057;
assign s[2039] = 8407081;
assign t[2039] = 2056;
assign s[2040] = 8405024;
assign t[2040] = 2055;
assign s[2041] = 8402969;
assign t[2041] = 2054;
assign s[2042] = 8400914;
assign t[2042] = 2053;
assign s[2043] = 8398861;
assign t[2043] = 2052;
assign s[2044] = 8396808;
assign t[2044] = 2051;
assign s[2045] = 8394757;
assign t[2045] = 2050;
assign s[2046] = 8392706;
assign t[2046] = 2049;
assign s[2047] = 8390657;
assign t[2047] = 2048;

wire [10:0] key;
assign key = bdata[22:12];

wire [11:0] A2;
assign A2 = bdata[11:0];

wire [24:0] S;
assign S = s[key];

wire [12:0] T;
assign T = t[key];

wire [24:0] S_TA_1;
assign S_TA_1 = (T * A2);

wire one;
assign one = !(|bdata[22:0]);

reg [24:0] S_TA_1_reg;
reg [24:0] S_reg;
reg one_reg_1;
reg s1_1;
reg [8:0] ea126_1;
reg [8:0] ea127_1;
reg [8:0] ea128_1;
reg [7:0] eb_1;
reg notzero_1;
reg flag1_1;
reg [4:0] address1_1;
reg [23:0] akasuu_1;

always@(posedge clk) begin
akasuu_1 <= {1'b1,adata[22:0]};
S_TA_1_reg <= S_TA_1;
S_reg <= S;
one_reg_1 <= one;
s1_1 <= adata[31] ^ bdata[31];
ea126_1 <= adata[30:23] + 126;
ea127_1 <= adata[30:23] + 127;
ea128_1 <= adata[30:23] + 128;
eb_1 <= bdata[30:23];
flag1_1 <= flag_in;
address1_1 <= address_in;
notzero_1 <= (|adata[30:23]);
end

wire [24:0] S_TA;
assign S_TA = S_reg - (S_TA_1_reg >> 12);

reg one_reg;
reg s1;
reg [8:0] ea126;
reg [8:0] ea127;
reg [8:0] ea128;
reg [7:0] eb;
reg [23:0] akasuu;
reg [23:0] bkasuu;
reg flag1;
reg [4:0] address1;
reg notzero_2;

always@(posedge clk) begin
akasuu <= akasuu_1;
bkasuu <= one_reg_1 ? S_TA[24:1] : S_TA[23:0];
one_reg <= one_reg_1;
s1 <= s1_1;
ea126 <= ea126_1;
ea127 <= ea127_1;
ea128 <= ea128_1;
eb <= eb_1;
flag1 <= flag1_1;
address1 <= address1_1;
notzero_2 <= notzero_1;
end

wire [13:0] a0;
assign a0 = akasuu[23:10];

wire [13:0] b0;
assign b0 = bkasuu[23:10];

wire [9:0] a1;
assign a1 = akasuu[9:0];

wire [9:0] b1;
assign b1 = bkasuu[9:0];

reg [27:0] a0b0;
reg [23:0] a1b0;
reg [23:0] a0b1;
reg [7:0] e;
reg [7:0] e_kuriage;
reg s2;
reg notzero;
reg flag2;
reg [4:0] address2;

always@(posedge clk) begin

a0b0 <= a0 * b0;

a1b0 <= a1 * b0;

a0b1 <= a0 * b1;

e <= one_reg ? ((ea127 < eb) ? 0 : ea127-eb) : ((ea126 < eb) ? 0 : ea126-eb);

e_kuriage <= one_reg ? ((ea127 < eb) ? 0 : ea128-eb) : ((ea126 < eb) ? 0 : ea127-eb);

s2 <= s1;

notzero <= notzero_2;

flag2 <= flag1;

address2 <= address1;


end

wire [14:0] a0b1tasua1b0;
assign a0b1tasua1b0 = a1b0[23:10] + a0b1[23:10] ;

wire [15:0] kekka_L;
assign kekka_L= a0b1tasua1b0 + a0b0[14:0];

wire [12:0] kekka_H_carry;
assign kekka_H_carry = a0b0[27:15] + 1;

wire [12:0] kekka_H_nocarry;
assign kekka_H_nocarry = a0b0[27:15];

wire carry;
assign carry = kekka_L[15];

wire [24:0] kekka;
assign kekka = carry ? {kekka_H_carry,kekka_L[14:3]} : {kekka_H_nocarry,kekka_L[14:3]};


wire [31:0] kotae;
assign kotae = notzero ? 
( kekka[24] ? {s2,e_kuriage,kekka[23:1]} : {s2,e,kekka[22:0]} ) : 0;

always@(posedge clk) begin
result <= kotae;
flag_out <= flag2;
address_out <= address2;
end
endmodule

`default_nettype wire
