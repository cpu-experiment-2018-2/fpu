module fdiv(
  input wire        en,
  input wire [31:0] adata,
  input wire [31:0] bdata,
  output reg [31:0] result,
  output reg        done,
  output reg        busy,
  input wire        clk,
  input wire        rstn
  );

//WAIT_ST
reg [31:0] wadata;
reg [31:0] wbdata;

//STAGE1
reg [31:0] adata1;
reg [31:0] bdata1;
reg [31:0] x02bai;
reg [31:0] x02jyou;

//STAGE2
reg [31:0] adata2;
reg [31:0] bdata2;
reg [31:0] x02bai2;
reg        ax02s1;
reg [8:0]  ax02e1;
reg [24:0] bdatakari;
reg [24:0] x2jyoukari;

//STAGE3
reg [31:0] adata3;
reg [31:0] bdata3;
reg [31:0] x02bai3;
reg [47:0] ax02jyoukekka;
reg        ax02jyous2;
reg [8:0]  ax02jyoue2;

//STAGE4
reg [31:0] adata4;
reg [31:0] bdata4;
reg [31:0] x02bai4;
reg [31:0] minusax02jyou;

//STAGE5
reg [31:0] adata5;
reg [31:0] bdata5;
reg        invbs1;
reg [7:0]  invbe1;
reg [24:0] invbdeka;
reg [24:0] invbchibi;
reg invbtashi1hiki0;

//STAGE6
reg [31:0] adata6;
reg [31:0] bdata6;
reg [24:0] invbkekka;
reg        invbs2;
reg [7:0]  invbe2;

//STAGE7
reg [31:0] adata7;
reg [31:0] bdata7;
reg [31:0] invb;

//STAGE8
reg        s1;
reg [8:0]  e1;
reg [24:0] adatakari;
reg [24:0] invbkari;
reg [8:0]  esyuuseia;
reg [8:0]  esyuuseib;

//STAGE9
reg [47:0] kekka;
reg        s2;
reg [8:0]  e2;
reg underflow;

typedef enum logic [3:0] {
  WAIT_ST,STAGE1,STAGE2,STAGE3,STAGE4,STAGE5,STAGE6,STAGE7,STAGE8,STAGE9
,STAGE10}state_type;
state_type state;

always@(posedge clk) begin
  if (~rstn) begin
    result <= 0;
    done   <= 0;
    busy   <= 0;
    state  <= WAIT_ST;
  end else if (state == WAIT_ST) begin
    done <= 0;
    if (en) begin
      state <= STAGE1;
      busy <= 1;
      wadata <= adata;
      wbdata <= bdata;
    end
  end else if (state == STAGE1) begin
    state <= STAGE2;
    adata1 <= wadata;
    bdata1 <= wbdata;

    if (wbdata[22:12] == 0) begin 
      x02bai <= 32'b00111111111111111111000000000010;
      x02jyou <= 32'b00111111011111111110000000000101;
    end else if (wbdata[22:12] == 1) begin 
      x02bai <= 32'b00111111111111111101000000001010;
      x02jyou <= 32'b00111111011111111010000000011101;
    end else if (wbdata[22:12] == 2) begin 
      x02bai <= 32'b00111111111111111011000000011010;
      x02jyou <= 32'b00111111011111110110000001001101;
    end else if (wbdata[22:12] == 3) begin 
      x02bai <= 32'b00111111111111111001000000110010;
      x02jyou <= 32'b00111111011111110010000010010101;
    end else if (wbdata[22:12] == 4) begin 
      x02bai <= 32'b00111111111111110111000001010010;
      x02jyou <= 32'b00111111011111101110000011110101;
    end else if (wbdata[22:12] == 5) begin 
      x02bai <= 32'b00111111111111110101000001111010;
      x02jyou <= 32'b00111111011111101010000101101100;
    end else if (wbdata[22:12] == 6) begin 
      x02bai <= 32'b00111111111111110011000010101001;
      x02jyou <= 32'b00111111011111100110000111111010;
    end else if (wbdata[22:12] == 7) begin 
      x02bai <= 32'b00111111111111110001000011100001;
      x02jyou <= 32'b00111111011111100010001010100001;
    end else if (wbdata[22:12] == 8) begin 
      x02bai <= 32'b00111111111111101111000100100001;
      x02jyou <= 32'b00111111011111011110001101100001;
    end else if (wbdata[22:12] == 9) begin 
      x02bai <= 32'b00111111111111101101000101101000;
      x02jyou <= 32'b00111111011111011010010000110110;
    end else if (wbdata[22:12] == 10) begin 
      x02bai <= 32'b00111111111111101011000110111000;
      x02jyou <= 32'b00111111011111010110010100100100;
    end else if (wbdata[22:12] == 11) begin 
      x02bai <= 32'b00111111111111101001001000001111;
      x02jyou <= 32'b00111111011111010010011000101001;
    end else if (wbdata[22:12] == 12) begin 
      x02bai <= 32'b00111111111111100111001001101110;
      x02jyou <= 32'b00111111011111001110011101000101;
    end else if (wbdata[22:12] == 13) begin 
      x02bai <= 32'b00111111111111100101001011010101;
      x02jyou <= 32'b00111111011111001010100001111001;
    end else if (wbdata[22:12] == 14) begin 
      x02bai <= 32'b00111111111111100011001101000100;
      x02jyou <= 32'b00111111011111000110100111000101;
    end else if (wbdata[22:12] == 15) begin 
      x02bai <= 32'b00111111111111100001001110111011;
      x02jyou <= 32'b00111111011111000010101100101001;
    end else if (wbdata[22:12] == 16) begin 
      x02bai <= 32'b00111111111111011111010000111001;
      x02jyou <= 32'b00111111011110111110110010100010;
    end else if (wbdata[22:12] == 17) begin 
      x02bai <= 32'b00111111111111011101010011000000;
      x02jyou <= 32'b00111111011110111010111000110100;
    end else if (wbdata[22:12] == 18) begin 
      x02bai <= 32'b00111111111111011011010101001110;
      x02jyou <= 32'b00111111011110110110111111011101;
    end else if (wbdata[22:12] == 19) begin 
      x02bai <= 32'b00111111111111011001010111100100;
      x02jyou <= 32'b00111111011110110011000110011100;
    end else if (wbdata[22:12] == 20) begin 
      x02bai <= 32'b00111111111111010111011010000001;
      x02jyou <= 32'b00111111011110101111001101110010;
    end else if (wbdata[22:12] == 21) begin 
      x02bai <= 32'b00111111111111010101011100100111;
      x02jyou <= 32'b00111111011110101011010101100001;
    end else if (wbdata[22:12] == 22) begin 
      x02bai <= 32'b00111111111111010011011111010100;
      x02jyou <= 32'b00111111011110100111011101100101;
    end else if (wbdata[22:12] == 23) begin 
      x02bai <= 32'b00111111111111010001100010001001;
      x02jyou <= 32'b00111111011110100011100110000001;
    end else if (wbdata[22:12] == 24) begin 
      x02bai <= 32'b00111111111111001111100101000110;
      x02jyou <= 32'b00111111011110011111101110110101;
    end else if (wbdata[22:12] == 25) begin 
      x02bai <= 32'b00111111111111001101101000001010;
      x02jyou <= 32'b00111111011110011011110111111101;
    end else if (wbdata[22:12] == 26) begin 
      x02bai <= 32'b00111111111111001011101011010110;
      x02jyou <= 32'b00111111011110011000000001011110;
    end else if (wbdata[22:12] == 27) begin 
      x02bai <= 32'b00111111111111001001101110101010;
      x02jyou <= 32'b00111111011110010100001011010101;
    end else if (wbdata[22:12] == 28) begin 
      x02bai <= 32'b00111111111111000111110010000101;
      x02jyou <= 32'b00111111011110010000010101100010;
    end else if (wbdata[22:12] == 29) begin 
      x02bai <= 32'b00111111111111000101110101101001;
      x02jyou <= 32'b00111111011110001100100000001001;
    end else if (wbdata[22:12] == 30) begin 
      x02bai <= 32'b00111111111111000011111001010011;
      x02jyou <= 32'b00111111011110001000101011000011;
    end else if (wbdata[22:12] == 31) begin 
      x02bai <= 32'b00111111111111000001111101000110;
      x02jyou <= 32'b00111111011110000100110110010110;
    end else if (wbdata[22:12] == 32) begin 
      x02bai <= 32'b00111111111111000000000001000000;
      x02jyou <= 32'b00111111011110000001000001111110;
    end else if (wbdata[22:12] == 33) begin 
      x02bai <= 32'b00111111111110111110000101000010;
      x02jyou <= 32'b00111111011101111101001101111110;
    end else if (wbdata[22:12] == 34) begin 
      x02bai <= 32'b00111111111110111100001001001011;
      x02jyou <= 32'b00111111011101111001011010010011;
    end else if (wbdata[22:12] == 35) begin 
      x02bai <= 32'b00111111111110111010001101011100;
      x02jyou <= 32'b00111111011101110101100110111111;
    end else if (wbdata[22:12] == 36) begin 
      x02bai <= 32'b00111111111110111000010001110101;
      x02jyou <= 32'b00111111011101110001110100000010;
    end else if (wbdata[22:12] == 37) begin 
      x02bai <= 32'b00111111111110110110010110010101;
      x02jyou <= 32'b00111111011101101110000001011010;
    end else if (wbdata[22:12] == 38) begin 
      x02bai <= 32'b00111111111110110100011010111101;
      x02jyou <= 32'b00111111011101101010001111001010;
    end else if (wbdata[22:12] == 39) begin 
      x02bai <= 32'b00111111111110110010011111101100;
      x02jyou <= 32'b00111111011101100110011101001111;
    end else if (wbdata[22:12] == 40) begin 
      x02bai <= 32'b00111111111110110000100100100011;
      x02jyou <= 32'b00111111011101100010101011101011;
    end else if (wbdata[22:12] == 41) begin 
      x02bai <= 32'b00111111111110101110101001100001;
      x02jyou <= 32'b00111111011101011110111010011100;
    end else if (wbdata[22:12] == 42) begin 
      x02bai <= 32'b00111111111110101100101110100111;
      x02jyou <= 32'b00111111011101011011001001100100;
    end else if (wbdata[22:12] == 43) begin 
      x02bai <= 32'b00111111111110101010110011110101;
      x02jyou <= 32'b00111111011101010111011001000011;
    end else if (wbdata[22:12] == 44) begin 
      x02bai <= 32'b00111111111110101000111001001001;
      x02jyou <= 32'b00111111011101010011101000110110;
    end else if (wbdata[22:12] == 45) begin 
      x02bai <= 32'b00111111111110100110111110100110;
      x02jyou <= 32'b00111111011101001111111001000001;
    end else if (wbdata[22:12] == 46) begin 
      x02bai <= 32'b00111111111110100101000100001010;
      x02jyou <= 32'b00111111011101001100001001100001;
    end else if (wbdata[22:12] == 47) begin 
      x02bai <= 32'b00111111111110100011001001110101;
      x02jyou <= 32'b00111111011101001000011010010110;
    end else if (wbdata[22:12] == 48) begin 
      x02bai <= 32'b00111111111110100001001111101000;
      x02jyou <= 32'b00111111011101000100101011100011;
    end else if (wbdata[22:12] == 49) begin 
      x02bai <= 32'b00111111111110011111010101100011;
      x02jyou <= 32'b00111111011101000000111101000110;
    end else if (wbdata[22:12] == 50) begin 
      x02bai <= 32'b00111111111110011101011011100100;
      x02jyou <= 32'b00111111011100111101001110111100;
    end else if (wbdata[22:12] == 51) begin 
      x02bai <= 32'b00111111111110011011100001101110;
      x02jyou <= 32'b00111111011100111001100001001011;
    end else if (wbdata[22:12] == 52) begin 
      x02bai <= 32'b00111111111110011001100111111110;
      x02jyou <= 32'b00111111011100110101110011101101;
    end else if (wbdata[22:12] == 53) begin 
      x02bai <= 32'b00111111111110010111101110010110;
      x02jyou <= 32'b00111111011100110010000110100101;
    end else if (wbdata[22:12] == 54) begin 
      x02bai <= 32'b00111111111110010101110100110110;
      x02jyou <= 32'b00111111011100101110011001110101;
    end else if (wbdata[22:12] == 55) begin 
      x02bai <= 32'b00111111111110010011111011011101;
      x02jyou <= 32'b00111111011100101010101101011001;
    end else if (wbdata[22:12] == 56) begin 
      x02bai <= 32'b00111111111110010010000010001011;
      x02jyou <= 32'b00111111011100100111000001010011;
    end else if (wbdata[22:12] == 57) begin 
      x02bai <= 32'b00111111111110010000001001000001;
      x02jyou <= 32'b00111111011100100011010101100010;
    end else if (wbdata[22:12] == 58) begin 
      x02bai <= 32'b00111111111110001110001111111110;
      x02jyou <= 32'b00111111011100011111101010000111;
    end else if (wbdata[22:12] == 59) begin 
      x02bai <= 32'b00111111111110001100010111000010;
      x02jyou <= 32'b00111111011100011011111111000001;
    end else if (wbdata[22:12] == 60) begin 
      x02bai <= 32'b00111111111110001010011110001110;
      x02jyou <= 32'b00111111011100011000010100010001;
    end else if (wbdata[22:12] == 61) begin 
      x02bai <= 32'b00111111111110001000100101100001;
      x02jyou <= 32'b00111111011100010100101001110110;
    end else if (wbdata[22:12] == 62) begin 
      x02bai <= 32'b00111111111110000110101100111011;
      x02jyou <= 32'b00111111011100010000111111101111;
    end else if (wbdata[22:12] == 63) begin 
      x02bai <= 32'b00111111111110000100110100011101;
      x02jyou <= 32'b00111111011100001101010101111111;
    end else if (wbdata[22:12] == 64) begin 
      x02bai <= 32'b00111111111110000010111100000110;
      x02jyou <= 32'b00111111011100001001101100100100;
    end else if (wbdata[22:12] == 65) begin 
      x02bai <= 32'b00111111111110000001000011110110;
      x02jyou <= 32'b00111111011100000110000011011110;
    end else if (wbdata[22:12] == 66) begin 
      x02bai <= 32'b00111111111101111111001011101110;
      x02jyou <= 32'b00111111011100000010011010101110;
    end else if (wbdata[22:12] == 67) begin 
      x02bai <= 32'b00111111111101111101010011101100;
      x02jyou <= 32'b00111111011011111110110010010000;
    end else if (wbdata[22:12] == 68) begin 
      x02bai <= 32'b00111111111101111011011011110010;
      x02jyou <= 32'b00111111011011111011001010001010;
    end else if (wbdata[22:12] == 69) begin 
      x02bai <= 32'b00111111111101111001100100000000;
      x02jyou <= 32'b00111111011011110111100010011001;
    end else if (wbdata[22:12] == 70) begin 
      x02bai <= 32'b00111111111101110111101100010100;
      x02jyou <= 32'b00111111011011110011111010111100;
    end else if (wbdata[22:12] == 71) begin 
      x02bai <= 32'b00111111111101110101110100110000;
      x02jyou <= 32'b00111111011011110000010011110101;
    end else if (wbdata[22:12] == 72) begin 
      x02bai <= 32'b00111111111101110011111101010011;
      x02jyou <= 32'b00111111011011101100101101000010;
    end else if (wbdata[22:12] == 73) begin 
      x02bai <= 32'b00111111111101110010000101111101;
      x02jyou <= 32'b00111111011011101001000110100100;
    end else if (wbdata[22:12] == 74) begin 
      x02bai <= 32'b00111111111101110000001110101111;
      x02jyou <= 32'b00111111011011100101100000011100;
    end else if (wbdata[22:12] == 75) begin 
      x02bai <= 32'b00111111111101101110010111100111;
      x02jyou <= 32'b00111111011011100001111010100110;
    end else if (wbdata[22:12] == 76) begin 
      x02bai <= 32'b00111111111101101100100000100111;
      x02jyou <= 32'b00111111011011011110010101000111;
    end else if (wbdata[22:12] == 77) begin 
      x02bai <= 32'b00111111111101101010101001101110;
      x02jyou <= 32'b00111111011011011010101111111101;
    end else if (wbdata[22:12] == 78) begin 
      x02bai <= 32'b00111111111101101000110010111100;
      x02jyou <= 32'b00111111011011010111001011000111;
    end else if (wbdata[22:12] == 79) begin 
      x02bai <= 32'b00111111111101100110111100010001;
      x02jyou <= 32'b00111111011011010011100110100101;
    end else if (wbdata[22:12] == 80) begin 
      x02bai <= 32'b00111111111101100101000101101110;
      x02jyou <= 32'b00111111011011010000000010011001;
    end else if (wbdata[22:12] == 81) begin 
      x02bai <= 32'b00111111111101100011001111010001;
      x02jyou <= 32'b00111111011011001100011110100000;
    end else if (wbdata[22:12] == 82) begin 
      x02bai <= 32'b00111111111101100001011000111100;
      x02jyou <= 32'b00111111011011001000111010111101;
    end else if (wbdata[22:12] == 83) begin 
      x02bai <= 32'b00111111111101011111100010101101;
      x02jyou <= 32'b00111111011011000101010111101101;
    end else if (wbdata[22:12] == 84) begin 
      x02bai <= 32'b00111111111101011101101100100110;
      x02jyou <= 32'b00111111011011000001110100110010;
    end else if (wbdata[22:12] == 85) begin 
      x02bai <= 32'b00111111111101011011110110100110;
      x02jyou <= 32'b00111111011010111110010010001100;
    end else if (wbdata[22:12] == 86) begin 
      x02bai <= 32'b00111111111101011010000000101101;
      x02jyou <= 32'b00111111011010111010101111111010;
    end else if (wbdata[22:12] == 87) begin 
      x02bai <= 32'b00111111111101011000001010111011;
      x02jyou <= 32'b00111111011010110111001101111101;
    end else if (wbdata[22:12] == 88) begin 
      x02bai <= 32'b00111111111101010110010101010000;
      x02jyou <= 32'b00111111011010110011101100010011;
    end else if (wbdata[22:12] == 89) begin 
      x02bai <= 32'b00111111111101010100011111101100;
      x02jyou <= 32'b00111111011010110000001010111110;
    end else if (wbdata[22:12] == 90) begin 
      x02bai <= 32'b00111111111101010010101010001111;
      x02jyou <= 32'b00111111011010101100101001111101;
    end else if (wbdata[22:12] == 91) begin 
      x02bai <= 32'b00111111111101010000110100111010;
      x02jyou <= 32'b00111111011010101001001001010010;
    end else if (wbdata[22:12] == 92) begin 
      x02bai <= 32'b00111111111101001110111111101011;
      x02jyou <= 32'b00111111011010100101101000111001;
    end else if (wbdata[22:12] == 93) begin 
      x02bai <= 32'b00111111111101001101001010100011;
      x02jyou <= 32'b00111111011010100010001000110100;
    end else if (wbdata[22:12] == 94) begin 
      x02bai <= 32'b00111111111101001011010101100010;
      x02jyou <= 32'b00111111011010011110101001000011;
    end else if (wbdata[22:12] == 95) begin 
      x02bai <= 32'b00111111111101001001100000101001;
      x02jyou <= 32'b00111111011010011011001001101001;
    end else if (wbdata[22:12] == 96) begin 
      x02bai <= 32'b00111111111101000111101011110110;
      x02jyou <= 32'b00111111011010010111101010100000;
    end else if (wbdata[22:12] == 97) begin 
      x02bai <= 32'b00111111111101000101110111001010;
      x02jyou <= 32'b00111111011010010100001011101011;
    end else if (wbdata[22:12] == 98) begin 
      x02bai <= 32'b00111111111101000100000010100101;
      x02jyou <= 32'b00111111011010010000101101001011;
    end else if (wbdata[22:12] == 99) begin 
      x02bai <= 32'b00111111111101000010001110000111;
      x02jyou <= 32'b00111111011010001101001110111110;
    end else if (wbdata[22:12] == 100) begin 
      x02bai <= 32'b00111111111101000000011001110000;
      x02jyou <= 32'b00111111011010001001110001000110;
    end else if (wbdata[22:12] == 101) begin 
      x02bai <= 32'b00111111111100111110100101100000;
      x02jyou <= 32'b00111111011010000110010011100001;
    end else if (wbdata[22:12] == 102) begin 
      x02bai <= 32'b00111111111100111100110001010111;
      x02jyou <= 32'b00111111011010000010110110010000;
    end else if (wbdata[22:12] == 103) begin 
      x02bai <= 32'b00111111111100111010111101010101;
      x02jyou <= 32'b00111111011001111111011001010011;
    end else if (wbdata[22:12] == 104) begin 
      x02bai <= 32'b00111111111100111001001001011001;
      x02jyou <= 32'b00111111011001111011111100101001;
    end else if (wbdata[22:12] == 105) begin 
      x02bai <= 32'b00111111111100110111010101100101;
      x02jyou <= 32'b00111111011001111000100000010100;
    end else if (wbdata[22:12] == 106) begin 
      x02bai <= 32'b00111111111100110101100001110111;
      x02jyou <= 32'b00111111011001110101000100010000;
    end else if (wbdata[22:12] == 107) begin 
      x02bai <= 32'b00111111111100110011101110010001;
      x02jyou <= 32'b00111111011001110001101000100011;
    end else if (wbdata[22:12] == 108) begin 
      x02bai <= 32'b00111111111100110001111010110001;
      x02jyou <= 32'b00111111011001101110001101001000;
    end else if (wbdata[22:12] == 109) begin 
      x02bai <= 32'b00111111111100110000000111011000;
      x02jyou <= 32'b00111111011001101010110010000000;
    end else if (wbdata[22:12] == 110) begin 
      x02bai <= 32'b00111111111100101110010100000110;
      x02jyou <= 32'b00111111011001100111010111001100;
    end else if (wbdata[22:12] == 111) begin 
      x02bai <= 32'b00111111111100101100100000111010;
      x02jyou <= 32'b00111111011001100011111100101010;
    end else if (wbdata[22:12] == 112) begin 
      x02bai <= 32'b00111111111100101010101101110110;
      x02jyou <= 32'b00111111011001100000100010011110;
    end else if (wbdata[22:12] == 113) begin 
      x02bai <= 32'b00111111111100101000111010111000;
      x02jyou <= 32'b00111111011001011101001000100011;
    end else if (wbdata[22:12] == 114) begin 
      x02bai <= 32'b00111111111100100111001000000001;
      x02jyou <= 32'b00111111011001011001101110111101;
    end else if (wbdata[22:12] == 115) begin 
      x02bai <= 32'b00111111111100100101010101010001;
      x02jyou <= 32'b00111111011001010110010101101010;
    end else if (wbdata[22:12] == 116) begin 
      x02bai <= 32'b00111111111100100011100010101000;
      x02jyou <= 32'b00111111011001010010111100101010;
    end else if (wbdata[22:12] == 117) begin 
      x02bai <= 32'b00111111111100100001110000000101;
      x02jyou <= 32'b00111111011001001111100011111101;
    end else if (wbdata[22:12] == 118) begin 
      x02bai <= 32'b00111111111100011111111101101010;
      x02jyou <= 32'b00111111011001001100001011100100;
    end else if (wbdata[22:12] == 119) begin 
      x02bai <= 32'b00111111111100011110001011010101;
      x02jyou <= 32'b00111111011001001000110011011110;
    end else if (wbdata[22:12] == 120) begin 
      x02bai <= 32'b00111111111100011100011001000110;
      x02jyou <= 32'b00111111011001000101011011101001;
    end else if (wbdata[22:12] == 121) begin 
      x02bai <= 32'b00111111111100011010100110111111;
      x02jyou <= 32'b00111111011001000010000100001010;
    end else if (wbdata[22:12] == 122) begin 
      x02bai <= 32'b00111111111100011000110100111110;
      x02jyou <= 32'b00111111011000111110101100111101;
    end else if (wbdata[22:12] == 123) begin 
      x02bai <= 32'b00111111111100010111000011000100;
      x02jyou <= 32'b00111111011000111011010110000011;
    end else if (wbdata[22:12] == 124) begin 
      x02bai <= 32'b00111111111100010101010001010001;
      x02jyou <= 32'b00111111011000110111111111011100;
    end else if (wbdata[22:12] == 125) begin 
      x02bai <= 32'b00111111111100010011011111100100;
      x02jyou <= 32'b00111111011000110100101001000111;
    end else if (wbdata[22:12] == 126) begin 
      x02bai <= 32'b00111111111100010001101101111110;
      x02jyou <= 32'b00111111011000110001010011000110;
    end else if (wbdata[22:12] == 127) begin 
      x02bai <= 32'b00111111111100001111111100011111;
      x02jyou <= 32'b00111111011000101101111101011000;
    end else if (wbdata[22:12] == 128) begin 
      x02bai <= 32'b00111111111100001110001011000110;
      x02jyou <= 32'b00111111011000101010100111111100;
    end else if (wbdata[22:12] == 129) begin 
      x02bai <= 32'b00111111111100001100011001110100;
      x02jyou <= 32'b00111111011000100111010010110011;
    end else if (wbdata[22:12] == 130) begin 
      x02bai <= 32'b00111111111100001010101000101001;
      x02jyou <= 32'b00111111011000100011111101111110;
    end else if (wbdata[22:12] == 131) begin 
      x02bai <= 32'b00111111111100001000110111100101;
      x02jyou <= 32'b00111111011000100000101001011100;
    end else if (wbdata[22:12] == 132) begin 
      x02bai <= 32'b00111111111100000111000110100111;
      x02jyou <= 32'b00111111011000011101010101001100;
    end else if (wbdata[22:12] == 133) begin 
      x02bai <= 32'b00111111111100000101010101101111;
      x02jyou <= 32'b00111111011000011010000001001101;
    end else if (wbdata[22:12] == 134) begin 
      x02bai <= 32'b00111111111100000011100100111110;
      x02jyou <= 32'b00111111011000010110101101100001;
    end else if (wbdata[22:12] == 135) begin 
      x02bai <= 32'b00111111111100000001110100010100;
      x02jyou <= 32'b00111111011000010011011010001001;
    end else if (wbdata[22:12] == 136) begin 
      x02bai <= 32'b00111111111100000000000011110001;
      x02jyou <= 32'b00111111011000010000000111000100;
    end else if (wbdata[22:12] == 137) begin 
      x02bai <= 32'b00111111111011111110010011010100;
      x02jyou <= 32'b00111111011000001100110100010000;
    end else if (wbdata[22:12] == 138) begin 
      x02bai <= 32'b00111111111011111100100010111110;
      x02jyou <= 32'b00111111011000001001100001110000;
    end else if (wbdata[22:12] == 139) begin 
      x02bai <= 32'b00111111111011111010110010101110;
      x02jyou <= 32'b00111111011000000110001111100001;
    end else if (wbdata[22:12] == 140) begin 
      x02bai <= 32'b00111111111011111001000010100101;
      x02jyou <= 32'b00111111011000000010111101100110;
    end else if (wbdata[22:12] == 141) begin 
      x02bai <= 32'b00111111111011110111010010100010;
      x02jyou <= 32'b00111111010111111111101011111100;
    end else if (wbdata[22:12] == 142) begin 
      x02bai <= 32'b00111111111011110101100010100110;
      x02jyou <= 32'b00111111010111111100011010100101;
    end else if (wbdata[22:12] == 143) begin 
      x02bai <= 32'b00111111111011110011110010110000;
      x02jyou <= 32'b00111111010111111001001001011111;
    end else if (wbdata[22:12] == 144) begin 
      x02bai <= 32'b00111111111011110010000011000001;
      x02jyou <= 32'b00111111010111110101111000101101;
    end else if (wbdata[22:12] == 145) begin 
      x02bai <= 32'b00111111111011110000010011011001;
      x02jyou <= 32'b00111111010111110010101000001101;
    end else if (wbdata[22:12] == 146) begin 
      x02bai <= 32'b00111111111011101110100011110111;
      x02jyou <= 32'b00111111010111101111010111111111;
    end else if (wbdata[22:12] == 147) begin 
      x02bai <= 32'b00111111111011101100110100011011;
      x02jyou <= 32'b00111111010111101100001000000011;
    end else if (wbdata[22:12] == 148) begin 
      x02bai <= 32'b00111111111011101011000101000110;
      x02jyou <= 32'b00111111010111101000111000011001;
    end else if (wbdata[22:12] == 149) begin 
      x02bai <= 32'b00111111111011101001010101111000;
      x02jyou <= 32'b00111111010111100101101001000010;
    end else if (wbdata[22:12] == 150) begin 
      x02bai <= 32'b00111111111011100111100110110000;
      x02jyou <= 32'b00111111010111100010011001111101;
    end else if (wbdata[22:12] == 151) begin 
      x02bai <= 32'b00111111111011100101110111101110;
      x02jyou <= 32'b00111111010111011111001011001001;
    end else if (wbdata[22:12] == 152) begin 
      x02bai <= 32'b00111111111011100100001000110011;
      x02jyou <= 32'b00111111010111011011111100101000;
    end else if (wbdata[22:12] == 153) begin 
      x02bai <= 32'b00111111111011100010011001111110;
      x02jyou <= 32'b00111111010111011000101110011000;
    end else if (wbdata[22:12] == 154) begin 
      x02bai <= 32'b00111111111011100000101011010000;
      x02jyou <= 32'b00111111010111010101100000011011;
    end else if (wbdata[22:12] == 155) begin 
      x02bai <= 32'b00111111111011011110111100101000;
      x02jyou <= 32'b00111111010111010010010010101111;
    end else if (wbdata[22:12] == 156) begin 
      x02bai <= 32'b00111111111011011101001110000111;
      x02jyou <= 32'b00111111010111001111000101010111;
    end else if (wbdata[22:12] == 157) begin 
      x02bai <= 32'b00111111111011011011011111101100;
      x02jyou <= 32'b00111111010111001011111000001111;
    end else if (wbdata[22:12] == 158) begin 
      x02bai <= 32'b00111111111011011001110001010111;
      x02jyou <= 32'b00111111010111001000101011011001;
    end else if (wbdata[22:12] == 159) begin 
      x02bai <= 32'b00111111111011011000000011001001;
      x02jyou <= 32'b00111111010111000101011110110101;
    end else if (wbdata[22:12] == 160) begin 
      x02bai <= 32'b00111111111011010110010101000001;
      x02jyou <= 32'b00111111010111000010010010100010;
    end else if (wbdata[22:12] == 161) begin 
      x02bai <= 32'b00111111111011010100100111000000;
      x02jyou <= 32'b00111111010110111111000110100011;
    end else if (wbdata[22:12] == 162) begin 
      x02bai <= 32'b00111111111011010010111001000101;
      x02jyou <= 32'b00111111010110111011111010110100;
    end else if (wbdata[22:12] == 163) begin 
      x02bai <= 32'b00111111111011010001001011010000;
      x02jyou <= 32'b00111111010110111000101111010111;
    end else if (wbdata[22:12] == 164) begin 
      x02bai <= 32'b00111111111011001111011101100010;
      x02jyou <= 32'b00111111010110110101100100001100;
    end else if (wbdata[22:12] == 165) begin 
      x02bai <= 32'b00111111111011001101101111111010;
      x02jyou <= 32'b00111111010110110010011001010010;
    end else if (wbdata[22:12] == 166) begin 
      x02bai <= 32'b00111111111011001100000010011000;
      x02jyou <= 32'b00111111010110101111001110101001;
    end else if (wbdata[22:12] == 167) begin 
      x02bai <= 32'b00111111111011001010010100111101;
      x02jyou <= 32'b00111111010110101100000100010011;
    end else if (wbdata[22:12] == 168) begin 
      x02bai <= 32'b00111111111011001000100111101000;
      x02jyou <= 32'b00111111010110101000111010001110;
    end else if (wbdata[22:12] == 169) begin 
      x02bai <= 32'b00111111111011000110111010011010;
      x02jyou <= 32'b00111111010110100101110000011100;
    end else if (wbdata[22:12] == 170) begin 
      x02bai <= 32'b00111111111011000101001101010001;
      x02jyou <= 32'b00111111010110100010100110111000;
    end else if (wbdata[22:12] == 171) begin 
      x02bai <= 32'b00111111111011000011100000001111;
      x02jyou <= 32'b00111111010110011111011101101000;
    end else if (wbdata[22:12] == 172) begin 
      x02bai <= 32'b00111111111011000001110011010011;
      x02jyou <= 32'b00111111010110011100010100101000;
    end else if (wbdata[22:12] == 173) begin 
      x02bai <= 32'b00111111111011000000000110011110;
      x02jyou <= 32'b00111111010110011001001011111011;
    end else if (wbdata[22:12] == 174) begin 
      x02bai <= 32'b00111111111010111110011001101111;
      x02jyou <= 32'b00111111010110010110000011011111;
    end else if (wbdata[22:12] == 175) begin 
      x02bai <= 32'b00111111111010111100101101000110;
      x02jyou <= 32'b00111111010110010010111011010100;
    end else if (wbdata[22:12] == 176) begin 
      x02bai <= 32'b00111111111010111011000000100011;
      x02jyou <= 32'b00111111010110001111110011011001;
    end else if (wbdata[22:12] == 177) begin 
      x02bai <= 32'b00111111111010111001010100000110;
      x02jyou <= 32'b00111111010110001100101011110000;
    end else if (wbdata[22:12] == 178) begin 
      x02bai <= 32'b00111111111010110111100111110000;
      x02jyou <= 32'b00111111010110001001100100011001;
    end else if (wbdata[22:12] == 179) begin 
      x02bai <= 32'b00111111111010110101111011100000;
      x02jyou <= 32'b00111111010110000110011101010010;
    end else if (wbdata[22:12] == 180) begin 
      x02bai <= 32'b00111111111010110100001111010110;
      x02jyou <= 32'b00111111010110000011010110011101;
    end else if (wbdata[22:12] == 181) begin 
      x02bai <= 32'b00111111111010110010100011010011;
      x02jyou <= 32'b00111111010110000000001111111010;
    end else if (wbdata[22:12] == 182) begin 
      x02bai <= 32'b00111111111010110000110111010101;
      x02jyou <= 32'b00111111010101111101001001100110;
    end else if (wbdata[22:12] == 183) begin 
      x02bai <= 32'b00111111111010101111001011011110;
      x02jyou <= 32'b00111111010101111010000011100100;
    end else if (wbdata[22:12] == 184) begin 
      x02bai <= 32'b00111111111010101101011111101101;
      x02jyou <= 32'b00111111010101110110111101110011;
    end else if (wbdata[22:12] == 185) begin 
      x02bai <= 32'b00111111111010101011110100000010;
      x02jyou <= 32'b00111111010101110011111000010011;
    end else if (wbdata[22:12] == 186) begin 
      x02bai <= 32'b00111111111010101010001000011110;
      x02jyou <= 32'b00111111010101110000110011000110;
    end else if (wbdata[22:12] == 187) begin 
      x02bai <= 32'b00111111111010101000011100111111;
      x02jyou <= 32'b00111111010101101101101110000111;
    end else if (wbdata[22:12] == 188) begin 
      x02bai <= 32'b00111111111010100110110001100111;
      x02jyou <= 32'b00111111010101101010101001011010;
    end else if (wbdata[22:12] == 189) begin 
      x02bai <= 32'b00111111111010100101000110010100;
      x02jyou <= 32'b00111111010101100111100100111101;
    end else if (wbdata[22:12] == 190) begin 
      x02bai <= 32'b00111111111010100011011011001000;
      x02jyou <= 32'b00111111010101100100100000110001;
    end else if (wbdata[22:12] == 191) begin 
      x02bai <= 32'b00111111111010100001110000000010;
      x02jyou <= 32'b00111111010101100001011100110111;
    end else if (wbdata[22:12] == 192) begin 
      x02bai <= 32'b00111111111010100000000101000011;
      x02jyou <= 32'b00111111010101011110011001001110;
    end else if (wbdata[22:12] == 193) begin 
      x02bai <= 32'b00111111111010011110011010001001;
      x02jyou <= 32'b00111111010101011011010101110101;
    end else if (wbdata[22:12] == 194) begin 
      x02bai <= 32'b00111111111010011100101111010101;
      x02jyou <= 32'b00111111010101011000010010101100;
    end else if (wbdata[22:12] == 195) begin 
      x02bai <= 32'b00111111111010011011000100101000;
      x02jyou <= 32'b00111111010101010101001111110101;
    end else if (wbdata[22:12] == 196) begin 
      x02bai <= 32'b00111111111010011001011010000000;
      x02jyou <= 32'b00111111010101010010001101001101;
    end else if (wbdata[22:12] == 197) begin 
      x02bai <= 32'b00111111111010010111101111011111;
      x02jyou <= 32'b00111111010101001111001010111000;
    end else if (wbdata[22:12] == 198) begin 
      x02bai <= 32'b00111111111010010110000101000011;
      x02jyou <= 32'b00111111010101001100001000110001;
    end else if (wbdata[22:12] == 199) begin 
      x02bai <= 32'b00111111111010010100011010101110;
      x02jyou <= 32'b00111111010101001001000110111100;
    end else if (wbdata[22:12] == 200) begin 
      x02bai <= 32'b00111111111010010010110000011111;
      x02jyou <= 32'b00111111010101000110000101011000;
    end else if (wbdata[22:12] == 201) begin 
      x02bai <= 32'b00111111111010010001000110010110;
      x02jyou <= 32'b00111111010101000011000100000100;
    end else if (wbdata[22:12] == 202) begin 
      x02bai <= 32'b00111111111010001111011100010011;
      x02jyou <= 32'b00111111010101000000000011000001;
    end else if (wbdata[22:12] == 203) begin 
      x02bai <= 32'b00111111111010001101110010010110;
      x02jyou <= 32'b00111111010100111101000010001110;
    end else if (wbdata[22:12] == 204) begin 
      x02bai <= 32'b00111111111010001100001000011111;
      x02jyou <= 32'b00111111010100111010000001101011;
    end else if (wbdata[22:12] == 205) begin 
      x02bai <= 32'b00111111111010001010011110101110;
      x02jyou <= 32'b00111111010100110111000001011001;
    end else if (wbdata[22:12] == 206) begin 
      x02bai <= 32'b00111111111010001000110101000011;
      x02jyou <= 32'b00111111010100110100000001010111;
    end else if (wbdata[22:12] == 207) begin 
      x02bai <= 32'b00111111111010000111001011011110;
      x02jyou <= 32'b00111111010100110001000001100110;
    end else if (wbdata[22:12] == 208) begin 
      x02bai <= 32'b00111111111010000101100001111110;
      x02jyou <= 32'b00111111010100101110000010000011;
    end else if (wbdata[22:12] == 209) begin 
      x02bai <= 32'b00111111111010000011111000100101;
      x02jyou <= 32'b00111111010100101011000010110010;
    end else if (wbdata[22:12] == 210) begin 
      x02bai <= 32'b00111111111010000010001111010010;
      x02jyou <= 32'b00111111010100101000000011110010;
    end else if (wbdata[22:12] == 211) begin 
      x02bai <= 32'b00111111111010000000100110000101;
      x02jyou <= 32'b00111111010100100101000101000001;
    end else if (wbdata[22:12] == 212) begin 
      x02bai <= 32'b00111111111001111110111100111110;
      x02jyou <= 32'b00111111010100100010000110100001;
    end else if (wbdata[22:12] == 213) begin 
      x02bai <= 32'b00111111111001111101010011111101;
      x02jyou <= 32'b00111111010100011111001000010010;
    end else if (wbdata[22:12] == 214) begin 
      x02bai <= 32'b00111111111001111011101011000001;
      x02jyou <= 32'b00111111010100011100001010010001;
    end else if (wbdata[22:12] == 215) begin 
      x02bai <= 32'b00111111111001111010000010001100;
      x02jyou <= 32'b00111111010100011001001100100001;
    end else if (wbdata[22:12] == 216) begin 
      x02bai <= 32'b00111111111001111000011001011101;
      x02jyou <= 32'b00111111010100010110001111000010;
    end else if (wbdata[22:12] == 217) begin 
      x02bai <= 32'b00111111111001110110110000110011;
      x02jyou <= 32'b00111111010100010011010001110010;
    end else if (wbdata[22:12] == 218) begin 
      x02bai <= 32'b00111111111001110101001000010000;
      x02jyou <= 32'b00111111010100010000010100110011;
    end else if (wbdata[22:12] == 219) begin 
      x02bai <= 32'b00111111111001110011011111110010;
      x02jyou <= 32'b00111111010100001101011000000011;
    end else if (wbdata[22:12] == 220) begin 
      x02bai <= 32'b00111111111001110001110111011010;
      x02jyou <= 32'b00111111010100001010011011100011;
    end else if (wbdata[22:12] == 221) begin 
      x02bai <= 32'b00111111111001110000001111001000;
      x02jyou <= 32'b00111111010100000111011111010011;
    end else if (wbdata[22:12] == 222) begin 
      x02bai <= 32'b00111111111001101110100110111100;
      x02jyou <= 32'b00111111010100000100100011010011;
    end else if (wbdata[22:12] == 223) begin 
      x02bai <= 32'b00111111111001101100111110110110;
      x02jyou <= 32'b00111111010100000001100111100100;
    end else if (wbdata[22:12] == 224) begin 
      x02bai <= 32'b00111111111001101011010110110110;
      x02jyou <= 32'b00111111010011111110101100000100;
    end else if (wbdata[22:12] == 225) begin 
      x02bai <= 32'b00111111111001101001101110111011;
      x02jyou <= 32'b00111111010011111011110000110011;
    end else if (wbdata[22:12] == 226) begin 
      x02bai <= 32'b00111111111001101000000111000111;
      x02jyou <= 32'b00111111010011111000110101110011;
    end else if (wbdata[22:12] == 227) begin 
      x02bai <= 32'b00111111111001100110011111011000;
      x02jyou <= 32'b00111111010011110101111011000010;
    end else if (wbdata[22:12] == 228) begin 
      x02bai <= 32'b00111111111001100100110111101111;
      x02jyou <= 32'b00111111010011110011000000100001;
    end else if (wbdata[22:12] == 229) begin 
      x02bai <= 32'b00111111111001100011010000001100;
      x02jyou <= 32'b00111111010011110000000110010000;
    end else if (wbdata[22:12] == 230) begin 
      x02bai <= 32'b00111111111001100001101000101110;
      x02jyou <= 32'b00111111010011101101001100001101;
    end else if (wbdata[22:12] == 231) begin 
      x02bai <= 32'b00111111111001100000000001010111;
      x02jyou <= 32'b00111111010011101010010010011100;
    end else if (wbdata[22:12] == 232) begin 
      x02bai <= 32'b00111111111001011110011010000101;
      x02jyou <= 32'b00111111010011100111011000111010;
    end else if (wbdata[22:12] == 233) begin 
      x02bai <= 32'b00111111111001011100110010111001;
      x02jyou <= 32'b00111111010011100100011111100111;
    end else if (wbdata[22:12] == 234) begin 
      x02bai <= 32'b00111111111001011011001011110011;
      x02jyou <= 32'b00111111010011100001100110100100;
    end else if (wbdata[22:12] == 235) begin 
      x02bai <= 32'b00111111111001011001100100110011;
      x02jyou <= 32'b00111111010011011110101101110001;
    end else if (wbdata[22:12] == 236) begin 
      x02bai <= 32'b00111111111001010111111101111000;
      x02jyou <= 32'b00111111010011011011110101001100;
    end else if (wbdata[22:12] == 237) begin 
      x02bai <= 32'b00111111111001010110010111000100;
      x02jyou <= 32'b00111111010011011000111100111001;
    end else if (wbdata[22:12] == 238) begin 
      x02bai <= 32'b00111111111001010100110000010101;
      x02jyou <= 32'b00111111010011010110000100110100;
    end else if (wbdata[22:12] == 239) begin 
      x02bai <= 32'b00111111111001010011001001101011;
      x02jyou <= 32'b00111111010011010011001100111101;
    end else if (wbdata[22:12] == 240) begin 
      x02bai <= 32'b00111111111001010001100011001000;
      x02jyou <= 32'b00111111010011010000010101011000;
    end else if (wbdata[22:12] == 241) begin 
      x02bai <= 32'b00111111111001001111111100101010;
      x02jyou <= 32'b00111111010011001101011110000001;
    end else if (wbdata[22:12] == 242) begin 
      x02bai <= 32'b00111111111001001110010110010010;
      x02jyou <= 32'b00111111010011001010100110111010;
    end else if (wbdata[22:12] == 243) begin 
      x02bai <= 32'b00111111111001001100110000000000;
      x02jyou <= 32'b00111111010011000111110000000011;
    end else if (wbdata[22:12] == 244) begin 
      x02bai <= 32'b00111111111001001011001001110011;
      x02jyou <= 32'b00111111010011000100111001011001;
    end else if (wbdata[22:12] == 245) begin 
      x02bai <= 32'b00111111111001001001100011101100;
      x02jyou <= 32'b00111111010011000010000011000000;
    end else if (wbdata[22:12] == 246) begin 
      x02bai <= 32'b00111111111001000111111101101011;
      x02jyou <= 32'b00111111010010111111001100110110;
    end else if (wbdata[22:12] == 247) begin 
      x02bai <= 32'b00111111111001000110010111101111;
      x02jyou <= 32'b00111111010010111100010110111010;
    end else if (wbdata[22:12] == 248) begin 
      x02bai <= 32'b00111111111001000100110001111001;
      x02jyou <= 32'b00111111010010111001100001001110;
    end else if (wbdata[22:12] == 249) begin 
      x02bai <= 32'b00111111111001000011001100001001;
      x02jyou <= 32'b00111111010010110110101011110010;
    end else if (wbdata[22:12] == 250) begin 
      x02bai <= 32'b00111111111001000001100110011111;
      x02jyou <= 32'b00111111010010110011110110100110;
    end else if (wbdata[22:12] == 251) begin 
      x02bai <= 32'b00111111111001000000000000111010;
      x02jyou <= 32'b00111111010010110001000001100111;
    end else if (wbdata[22:12] == 252) begin 
      x02bai <= 32'b00111111111000111110011011011010;
      x02jyou <= 32'b00111111010010101110001100110111;
    end else if (wbdata[22:12] == 253) begin 
      x02bai <= 32'b00111111111000111100110110000001;
      x02jyou <= 32'b00111111010010101011011000011000;
    end else if (wbdata[22:12] == 254) begin 
      x02bai <= 32'b00111111111000111011010000101101;
      x02jyou <= 32'b00111111010010101000100100000111;
    end else if (wbdata[22:12] == 255) begin 
      x02bai <= 32'b00111111111000111001101011011111;
      x02jyou <= 32'b00111111010010100101110000000101;
    end else if (wbdata[22:12] == 256) begin 
      x02bai <= 32'b00111111111000111000000110010110;
      x02jyou <= 32'b00111111010010100010111100010010;
    end else if (wbdata[22:12] == 257) begin 
      x02bai <= 32'b00111111111000110110100001010011;
      x02jyou <= 32'b00111111010010100000001000101110;
    end else if (wbdata[22:12] == 258) begin 
      x02bai <= 32'b00111111111000110100111100010101;
      x02jyou <= 32'b00111111010010011101010101011000;
    end else if (wbdata[22:12] == 259) begin 
      x02bai <= 32'b00111111111000110011010111011110;
      x02jyou <= 32'b00111111010010011010100010010011;
    end else if (wbdata[22:12] == 260) begin 
      x02bai <= 32'b00111111111000110001110010101011;
      x02jyou <= 32'b00111111010010010111101111011010;
    end else if (wbdata[22:12] == 261) begin 
      x02bai <= 32'b00111111111000110000001101111111;
      x02jyou <= 32'b00111111010010010100111100110011;
    end else if (wbdata[22:12] == 262) begin 
      x02bai <= 32'b00111111111000101110101001010111;
      x02jyou <= 32'b00111111010010010010001010011000;
    end else if (wbdata[22:12] == 263) begin 
      x02bai <= 32'b00111111111000101101000100110110;
      x02jyou <= 32'b00111111010010001111011000001110;
    end else if (wbdata[22:12] == 264) begin 
      x02bai <= 32'b00111111111000101011100000011010;
      x02jyou <= 32'b00111111010010001100100110010010;
    end else if (wbdata[22:12] == 265) begin 
      x02bai <= 32'b00111111111000101001111100000100;
      x02jyou <= 32'b00111111010010001001110100100110;
    end else if (wbdata[22:12] == 266) begin 
      x02bai <= 32'b00111111111000101000010111110011;
      x02jyou <= 32'b00111111010010000111000011000111;
    end else if (wbdata[22:12] == 267) begin 
      x02bai <= 32'b00111111111000100110110011100111;
      x02jyou <= 32'b00111111010010000100010001110110;
    end else if (wbdata[22:12] == 268) begin 
      x02bai <= 32'b00111111111000100101001111100010;
      x02jyou <= 32'b00111111010010000001100000110111;
    end else if (wbdata[22:12] == 269) begin 
      x02bai <= 32'b00111111111000100011101011100001;
      x02jyou <= 32'b00111111010001111110110000000011;
    end else if (wbdata[22:12] == 270) begin 
      x02bai <= 32'b00111111111000100010000111100111;
      x02jyou <= 32'b00111111010001111011111111100000;
    end else if (wbdata[22:12] == 271) begin 
      x02bai <= 32'b00111111111000100000100011110001;
      x02jyou <= 32'b00111111010001111001001111001010;
    end else if (wbdata[22:12] == 272) begin 
      x02bai <= 32'b00111111111000011111000000000010;
      x02jyou <= 32'b00111111010001110110011111000101;
    end else if (wbdata[22:12] == 273) begin 
      x02bai <= 32'b00111111111000011101011100010111;
      x02jyou <= 32'b00111111010001110011101111001011;
    end else if (wbdata[22:12] == 274) begin 
      x02bai <= 32'b00111111111000011011111000110011;
      x02jyou <= 32'b00111111010001110000111111100011;
    end else if (wbdata[22:12] == 275) begin 
      x02bai <= 32'b00111111111000011010010101010011;
      x02jyou <= 32'b00111111010001101110010000000111;
    end else if (wbdata[22:12] == 276) begin 
      x02bai <= 32'b00111111111000011000110001111010;
      x02jyou <= 32'b00111111010001101011100000111100;
    end else if (wbdata[22:12] == 277) begin 
      x02bai <= 32'b00111111111000010111001110100101;
      x02jyou <= 32'b00111111010001101000110001111100;
    end else if (wbdata[22:12] == 278) begin 
      x02bai <= 32'b00111111111000010101101011010110;
      x02jyou <= 32'b00111111010001100110000011001100;
    end else if (wbdata[22:12] == 279) begin 
      x02bai <= 32'b00111111111000010100001000001101;
      x02jyou <= 32'b00111111010001100011010100101100;
    end else if (wbdata[22:12] == 280) begin 
      x02bai <= 32'b00111111111000010010100101001001;
      x02jyou <= 32'b00111111010001100000100110011001;
    end else if (wbdata[22:12] == 281) begin 
      x02bai <= 32'b00111111111000010001000010001011;
      x02jyou <= 32'b00111111010001011101111000010101;
    end else if (wbdata[22:12] == 282) begin 
      x02bai <= 32'b00111111111000001111011111010010;
      x02jyou <= 32'b00111111010001011011001010011111;
    end else if (wbdata[22:12] == 283) begin 
      x02bai <= 32'b00111111111000001101111100011110;
      x02jyou <= 32'b00111111010001011000011100110111;
    end else if (wbdata[22:12] == 284) begin 
      x02bai <= 32'b00111111111000001100011001110000;
      x02jyou <= 32'b00111111010001010101101111011110;
    end else if (wbdata[22:12] == 285) begin 
      x02bai <= 32'b00111111111000001010110111000111;
      x02jyou <= 32'b00111111010001010011000010010010;
    end else if (wbdata[22:12] == 286) begin 
      x02bai <= 32'b00111111111000001001010100100100;
      x02jyou <= 32'b00111111010001010000010101010110;
    end else if (wbdata[22:12] == 287) begin 
      x02bai <= 32'b00111111111000000111110010000110;
      x02jyou <= 32'b00111111010001001101101000100111;
    end else if (wbdata[22:12] == 288) begin 
      x02bai <= 32'b00111111111000000110001111101101;
      x02jyou <= 32'b00111111010001001010111100000110;
    end else if (wbdata[22:12] == 289) begin 
      x02bai <= 32'b00111111111000000100101101011010;
      x02jyou <= 32'b00111111010001001000001111110100;
    end else if (wbdata[22:12] == 290) begin 
      x02bai <= 32'b00111111111000000011001011001100;
      x02jyou <= 32'b00111111010001000101100011101111;
    end else if (wbdata[22:12] == 291) begin 
      x02bai <= 32'b00111111111000000001101001000100;
      x02jyou <= 32'b00111111010001000010110111111010;
    end else if (wbdata[22:12] == 292) begin 
      x02bai <= 32'b00111111111000000000000111000001;
      x02jyou <= 32'b00111111010001000000001100010010;
    end else if (wbdata[22:12] == 293) begin 
      x02bai <= 32'b00111111110111111110100101000011;
      x02jyou <= 32'b00111111010000111101100000110111;
    end else if (wbdata[22:12] == 294) begin 
      x02bai <= 32'b00111111110111111101000011001011;
      x02jyou <= 32'b00111111010000111010110101101100;
    end else if (wbdata[22:12] == 295) begin 
      x02bai <= 32'b00111111110111111011100001011000;
      x02jyou <= 32'b00111111010000111000001010101110;
    end else if (wbdata[22:12] == 296) begin 
      x02bai <= 32'b00111111110111111001111111101010;
      x02jyou <= 32'b00111111010000110101011111111110;
    end else if (wbdata[22:12] == 297) begin 
      x02bai <= 32'b00111111110111111000011110000010;
      x02jyou <= 32'b00111111010000110010110101011100;
    end else if (wbdata[22:12] == 298) begin 
      x02bai <= 32'b00111111110111110110111100011111;
      x02jyou <= 32'b00111111010000110000001011001000;
    end else if (wbdata[22:12] == 299) begin 
      x02bai <= 32'b00111111110111110101011011000001;
      x02jyou <= 32'b00111111010000101101100001000010;
    end else if (wbdata[22:12] == 300) begin 
      x02bai <= 32'b00111111110111110011111001101001;
      x02jyou <= 32'b00111111010000101010110111001010;
    end else if (wbdata[22:12] == 301) begin 
      x02bai <= 32'b00111111110111110010011000010101;
      x02jyou <= 32'b00111111010000101000001101011110;
    end else if (wbdata[22:12] == 302) begin 
      x02bai <= 32'b00111111110111110000110111001000;
      x02jyou <= 32'b00111111010000100101100100000011;
    end else if (wbdata[22:12] == 303) begin 
      x02bai <= 32'b00111111110111101111010101111111;
      x02jyou <= 32'b00111111010000100010111010110100;
    end else if (wbdata[22:12] == 304) begin 
      x02bai <= 32'b00111111110111101101110100111100;
      x02jyou <= 32'b00111111010000100000010001110011;
    end else if (wbdata[22:12] == 305) begin 
      x02bai <= 32'b00111111110111101100010011111110;
      x02jyou <= 32'b00111111010000011101101001000000;
    end else if (wbdata[22:12] == 306) begin 
      x02bai <= 32'b00111111110111101010110011000101;
      x02jyou <= 32'b00111111010000011011000000011010;
    end else if (wbdata[22:12] == 307) begin 
      x02bai <= 32'b00111111110111101001010010010010;
      x02jyou <= 32'b00111111010000011000011000000011;
    end else if (wbdata[22:12] == 308) begin 
      x02bai <= 32'b00111111110111100111110001100100;
      x02jyou <= 32'b00111111010000010101101111111010;
    end else if (wbdata[22:12] == 309) begin 
      x02bai <= 32'b00111111110111100110010000111011;
      x02jyou <= 32'b00111111010000010011000111111110;
    end else if (wbdata[22:12] == 310) begin 
      x02bai <= 32'b00111111110111100100110000010111;
      x02jyou <= 32'b00111111010000010000100000001111;
    end else if (wbdata[22:12] == 311) begin 
      x02bai <= 32'b00111111110111100011001111111001;
      x02jyou <= 32'b00111111010000001101111000101110;
    end else if (wbdata[22:12] == 312) begin 
      x02bai <= 32'b00111111110111100001101111100000;
      x02jyou <= 32'b00111111010000001011010001011100;
    end else if (wbdata[22:12] == 313) begin 
      x02bai <= 32'b00111111110111100000001111001100;
      x02jyou <= 32'b00111111010000001000101010010110;
    end else if (wbdata[22:12] == 314) begin 
      x02bai <= 32'b00111111110111011110101110111101;
      x02jyou <= 32'b00111111010000000110000011011101;
    end else if (wbdata[22:12] == 315) begin 
      x02bai <= 32'b00111111110111011101001110110100;
      x02jyou <= 32'b00111111010000000011011100110100;
    end else if (wbdata[22:12] == 316) begin 
      x02bai <= 32'b00111111110111011011101110101111;
      x02jyou <= 32'b00111111010000000000110110010110;
    end else if (wbdata[22:12] == 317) begin 
      x02bai <= 32'b00111111110111011010001110110000;
      x02jyou <= 32'b00111111001111111110010000000111;
    end else if (wbdata[22:12] == 318) begin 
      x02bai <= 32'b00111111110111011000101110110110;
      x02jyou <= 32'b00111111001111111011101010000100;
    end else if (wbdata[22:12] == 319) begin 
      x02bai <= 32'b00111111110111010111001111000010;
      x02jyou <= 32'b00111111001111111001000100010001;
    end else if (wbdata[22:12] == 320) begin 
      x02bai <= 32'b00111111110111010101101111010010;
      x02jyou <= 32'b00111111001111110110011110101010;
    end else if (wbdata[22:12] == 321) begin 
      x02bai <= 32'b00111111110111010100001111101000;
      x02jyou <= 32'b00111111001111110011111001010001;
    end else if (wbdata[22:12] == 322) begin 
      x02bai <= 32'b00111111110111010010110000000011;
      x02jyou <= 32'b00111111001111110001010100000101;
    end else if (wbdata[22:12] == 323) begin 
      x02bai <= 32'b00111111110111010001010000100011;
      x02jyou <= 32'b00111111001111101110101111000110;
    end else if (wbdata[22:12] == 324) begin 
      x02bai <= 32'b00111111110111001111110001001000;
      x02jyou <= 32'b00111111001111101100001010010100;
    end else if (wbdata[22:12] == 325) begin 
      x02bai <= 32'b00111111110111001110010001110010;
      x02jyou <= 32'b00111111001111101001100101110000;
    end else if (wbdata[22:12] == 326) begin 
      x02bai <= 32'b00111111110111001100110010100001;
      x02jyou <= 32'b00111111001111100111000001011000;
    end else if (wbdata[22:12] == 327) begin 
      x02bai <= 32'b00111111110111001011010011010110;
      x02jyou <= 32'b00111111001111100100011101010000;
    end else if (wbdata[22:12] == 328) begin 
      x02bai <= 32'b00111111110111001001110100001111;
      x02jyou <= 32'b00111111001111100001111001010010;
    end else if (wbdata[22:12] == 329) begin 
      x02bai <= 32'b00111111110111001000010101001110;
      x02jyou <= 32'b00111111001111011111010101100011;
    end else if (wbdata[22:12] == 330) begin 
      x02bai <= 32'b00111111110111000110110110010010;
      x02jyou <= 32'b00111111001111011100110010000010;
    end else if (wbdata[22:12] == 331) begin 
      x02bai <= 32'b00111111110111000101010111011011;
      x02jyou <= 32'b00111111001111011010001110101101;
    end else if (wbdata[22:12] == 332) begin 
      x02bai <= 32'b00111111110111000011111000101001;
      x02jyou <= 32'b00111111001111010111101011100110;
    end else if (wbdata[22:12] == 333) begin 
      x02bai <= 32'b00111111110111000010011001111100;
      x02jyou <= 32'b00111111001111010101001000101011;
    end else if (wbdata[22:12] == 334) begin 
      x02bai <= 32'b00111111110111000000111011010101;
      x02jyou <= 32'b00111111001111010010100101111111;
    end else if (wbdata[22:12] == 335) begin 
      x02bai <= 32'b00111111110110111111011100110010;
      x02jyou <= 32'b00111111001111010000000011011110;
    end else if (wbdata[22:12] == 336) begin 
      x02bai <= 32'b00111111110110111101111110010100;
      x02jyou <= 32'b00111111001111001101100001001010;
    end else if (wbdata[22:12] == 337) begin 
      x02bai <= 32'b00111111110110111100011111111100;
      x02jyou <= 32'b00111111001111001010111111000101;
    end else if (wbdata[22:12] == 338) begin 
      x02bai <= 32'b00111111110110111011000001101000;
      x02jyou <= 32'b00111111001111001000011101001011;
    end else if (wbdata[22:12] == 339) begin 
      x02bai <= 32'b00111111110110111001100011011010;
      x02jyou <= 32'b00111111001111000101111011100000;
    end else if (wbdata[22:12] == 340) begin 
      x02bai <= 32'b00111111110110111000000101010001;
      x02jyou <= 32'b00111111001111000011011010000010;
    end else if (wbdata[22:12] == 341) begin 
      x02bai <= 32'b00111111110110110110100111001100;
      x02jyou <= 32'b00111111001111000000111000101111;
    end else if (wbdata[22:12] == 342) begin 
      x02bai <= 32'b00111111110110110101001001001101;
      x02jyou <= 32'b00111111001110111110010111101010;
    end else if (wbdata[22:12] == 343) begin 
      x02bai <= 32'b00111111110110110011101011010011;
      x02jyou <= 32'b00111111001110111011110110110011;
    end else if (wbdata[22:12] == 344) begin 
      x02bai <= 32'b00111111110110110010001101011110;
      x02jyou <= 32'b00111111001110111001010110001000;
    end else if (wbdata[22:12] == 345) begin 
      x02bai <= 32'b00111111110110110000101111101110;
      x02jyou <= 32'b00111111001110110110110101101010;
    end else if (wbdata[22:12] == 346) begin 
      x02bai <= 32'b00111111110110101111010010000010;
      x02jyou <= 32'b00111111001110110100010101010111;
    end else if (wbdata[22:12] == 347) begin 
      x02bai <= 32'b00111111110110101101110100011100;
      x02jyou <= 32'b00111111001110110001110101010011;
    end else if (wbdata[22:12] == 348) begin 
      x02bai <= 32'b00111111110110101100010110111011;
      x02jyou <= 32'b00111111001110101111010101011011;
    end else if (wbdata[22:12] == 349) begin 
      x02bai <= 32'b00111111110110101010111001011111;
      x02jyou <= 32'b00111111001110101100110101110001;
    end else if (wbdata[22:12] == 350) begin 
      x02bai <= 32'b00111111110110101001011100001000;
      x02jyou <= 32'b00111111001110101010010110010011;
    end else if (wbdata[22:12] == 351) begin 
      x02bai <= 32'b00111111110110100111111110110110;
      x02jyou <= 32'b00111111001110100111110111000010;
    end else if (wbdata[22:12] == 352) begin 
      x02bai <= 32'b00111111110110100110100001101000;
      x02jyou <= 32'b00111111001110100101010111111100;
    end else if (wbdata[22:12] == 353) begin 
      x02bai <= 32'b00111111110110100101000100100000;
      x02jyou <= 32'b00111111001110100010111001000100;
    end else if (wbdata[22:12] == 354) begin 
      x02bai <= 32'b00111111110110100011100111011101;
      x02jyou <= 32'b00111111001110100000011010011001;
    end else if (wbdata[22:12] == 355) begin 
      x02bai <= 32'b00111111110110100010001010011110;
      x02jyou <= 32'b00111111001110011101111011111010;
    end else if (wbdata[22:12] == 356) begin 
      x02bai <= 32'b00111111110110100000101101100101;
      x02jyou <= 32'b00111111001110011011011101101001;
    end else if (wbdata[22:12] == 357) begin 
      x02bai <= 32'b00111111110110011111010000110001;
      x02jyou <= 32'b00111111001110011000111111100100;
    end else if (wbdata[22:12] == 358) begin 
      x02bai <= 32'b00111111110110011101110100000001;
      x02jyou <= 32'b00111111001110010110100001101010;
    end else if (wbdata[22:12] == 359) begin 
      x02bai <= 32'b00111111110110011100010111010110;
      x02jyou <= 32'b00111111001110010100000011111110;
    end else if (wbdata[22:12] == 360) begin 
      x02bai <= 32'b00111111110110011010111010110001;
      x02jyou <= 32'b00111111001110010001100110011111;
    end else if (wbdata[22:12] == 361) begin 
      x02bai <= 32'b00111111110110011001011110010000;
      x02jyou <= 32'b00111111001110001111001001001100;
    end else if (wbdata[22:12] == 362) begin 
      x02bai <= 32'b00111111110110011000000001110100;
      x02jyou <= 32'b00111111001110001100101100000101;
    end else if (wbdata[22:12] == 363) begin 
      x02bai <= 32'b00111111110110010110100101011101;
      x02jyou <= 32'b00111111001110001010001111001011;
    end else if (wbdata[22:12] == 364) begin 
      x02bai <= 32'b00111111110110010101001001001011;
      x02jyou <= 32'b00111111001110000111110010011110;
    end else if (wbdata[22:12] == 365) begin 
      x02bai <= 32'b00111111110110010011101100111110;
      x02jyou <= 32'b00111111001110000101010101111101;
    end else if (wbdata[22:12] == 366) begin 
      x02bai <= 32'b00111111110110010010010000110110;
      x02jyou <= 32'b00111111001110000010111001101001;
    end else if (wbdata[22:12] == 367) begin 
      x02bai <= 32'b00111111110110010000110100110010;
      x02jyou <= 32'b00111111001110000000011101011111;
    end else if (wbdata[22:12] == 368) begin 
      x02bai <= 32'b00111111110110001111011000110100;
      x02jyou <= 32'b00111111001101111110000001100101;
    end else if (wbdata[22:12] == 369) begin 
      x02bai <= 32'b00111111110110001101111100111010;
      x02jyou <= 32'b00111111001101111011100101110101;
    end else if (wbdata[22:12] == 370) begin 
      x02bai <= 32'b00111111110110001100100001000110;
      x02jyou <= 32'b00111111001101111001001010010011;
    end else if (wbdata[22:12] == 371) begin 
      x02bai <= 32'b00111111110110001011000101010110;
      x02jyou <= 32'b00111111001101110110101110111100;
    end else if (wbdata[22:12] == 372) begin 
      x02bai <= 32'b00111111110110001001101001101011;
      x02jyou <= 32'b00111111001101110100010011110010;
    end else if (wbdata[22:12] == 373) begin 
      x02bai <= 32'b00111111110110001000001110000100;
      x02jyou <= 32'b00111111001101110001111000110010;
    end else if (wbdata[22:12] == 374) begin 
      x02bai <= 32'b00111111110110000110110010100011;
      x02jyou <= 32'b00111111001101101111011110000001;
    end else if (wbdata[22:12] == 375) begin 
      x02bai <= 32'b00111111110110000101010111000111;
      x02jyou <= 32'b00111111001101101101000011011101;
    end else if (wbdata[22:12] == 376) begin 
      x02bai <= 32'b00111111110110000011111011101111;
      x02jyou <= 32'b00111111001101101010101001000011;
    end else if (wbdata[22:12] == 377) begin 
      x02bai <= 32'b00111111110110000010100000011100;
      x02jyou <= 32'b00111111001101101000001110110110;
    end else if (wbdata[22:12] == 378) begin 
      x02bai <= 32'b00111111110110000001000101001110;
      x02jyou <= 32'b00111111001101100101110100110101;
    end else if (wbdata[22:12] == 379) begin 
      x02bai <= 32'b00111111110101111111101010000101;
      x02jyou <= 32'b00111111001101100011011011000001;
    end else if (wbdata[22:12] == 380) begin 
      x02bai <= 32'b00111111110101111110001111000000;
      x02jyou <= 32'b00111111001101100001000001010111;
    end else if (wbdata[22:12] == 381) begin 
      x02bai <= 32'b00111111110101111100110100000001;
      x02jyou <= 32'b00111111001101011110100111111100;
    end else if (wbdata[22:12] == 382) begin 
      x02bai <= 32'b00111111110101111011011001000110;
      x02jyou <= 32'b00111111001101011100001110101011;
    end else if (wbdata[22:12] == 383) begin 
      x02bai <= 32'b00111111110101111001111110010000;
      x02jyou <= 32'b00111111001101011001110101100111;
    end else if (wbdata[22:12] == 384) begin 
      x02bai <= 32'b00111111110101111000100011011110;
      x02jyou <= 32'b00111111001101010111011100101110;
    end else if (wbdata[22:12] == 385) begin 
      x02bai <= 32'b00111111110101110111001000110010;
      x02jyou <= 32'b00111111001101010101000100000011;
    end else if (wbdata[22:12] == 386) begin 
      x02bai <= 32'b00111111110101110101101110001010;
      x02jyou <= 32'b00111111001101010010101011100011;
    end else if (wbdata[22:12] == 387) begin 
      x02bai <= 32'b00111111110101110100010011100111;
      x02jyou <= 32'b00111111001101010000010011001111;
    end else if (wbdata[22:12] == 388) begin 
      x02bai <= 32'b00111111110101110010111001001001;
      x02jyou <= 32'b00111111001101001101111011000111;
    end else if (wbdata[22:12] == 389) begin 
      x02bai <= 32'b00111111110101110001011110110000;
      x02jyou <= 32'b00111111001101001011100011001100;
    end else if (wbdata[22:12] == 390) begin 
      x02bai <= 32'b00111111110101110000000100011011;
      x02jyou <= 32'b00111111001101001001001011011011;
    end else if (wbdata[22:12] == 391) begin 
      x02bai <= 32'b00111111110101101110101010001011;
      x02jyou <= 32'b00111111001101000110110011110111;
    end else if (wbdata[22:12] == 392) begin 
      x02bai <= 32'b00111111110101101101010000000000;
      x02jyou <= 32'b00111111001101000100011100100000;
    end else if (wbdata[22:12] == 393) begin 
      x02bai <= 32'b00111111110101101011110101111001;
      x02jyou <= 32'b00111111001101000010000101010011;
    end else if (wbdata[22:12] == 394) begin 
      x02bai <= 32'b00111111110101101010011011110111;
      x02jyou <= 32'b00111111001100111111101110010010;
    end else if (wbdata[22:12] == 395) begin 
      x02bai <= 32'b00111111110101101001000001111010;
      x02jyou <= 32'b00111111001100111101010111011110;
    end else if (wbdata[22:12] == 396) begin 
      x02bai <= 32'b00111111110101100111101000000010;
      x02jyou <= 32'b00111111001100111011000000110101;
    end else if (wbdata[22:12] == 397) begin 
      x02bai <= 32'b00111111110101100110001110001110;
      x02jyou <= 32'b00111111001100111000101010011000;
    end else if (wbdata[22:12] == 398) begin 
      x02bai <= 32'b00111111110101100100110100011111;
      x02jyou <= 32'b00111111001100110110010100000111;
    end else if (wbdata[22:12] == 399) begin 
      x02bai <= 32'b00111111110101100011011010110101;
      x02jyou <= 32'b00111111001100110011111110000010;
    end else if (wbdata[22:12] == 400) begin 
      x02bai <= 32'b00111111110101100010000001001111;
      x02jyou <= 32'b00111111001100110001101000001000;
    end else if (wbdata[22:12] == 401) begin 
      x02bai <= 32'b00111111110101100000100111101110;
      x02jyou <= 32'b00111111001100101111010010011010;
    end else if (wbdata[22:12] == 402) begin 
      x02bai <= 32'b00111111110101011111001110010010;
      x02jyou <= 32'b00111111001100101100111100111001;
    end else if (wbdata[22:12] == 403) begin 
      x02bai <= 32'b00111111110101011101110100111010;
      x02jyou <= 32'b00111111001100101010100111100010;
    end else if (wbdata[22:12] == 404) begin 
      x02bai <= 32'b00111111110101011100011011101000;
      x02jyou <= 32'b00111111001100101000010010011001;
    end else if (wbdata[22:12] == 405) begin 
      x02bai <= 32'b00111111110101011011000010011001;
      x02jyou <= 32'b00111111001100100101111101011000;
    end else if (wbdata[22:12] == 406) begin 
      x02bai <= 32'b00111111110101011001101001010000;
      x02jyou <= 32'b00111111001100100011101000100110;
    end else if (wbdata[22:12] == 407) begin 
      x02bai <= 32'b00111111110101011000010000001011;
      x02jyou <= 32'b00111111001100100001010011111110;
    end else if (wbdata[22:12] == 408) begin 
      x02bai <= 32'b00111111110101010110110111001010;
      x02jyou <= 32'b00111111001100011110111111100001;
    end else if (wbdata[22:12] == 409) begin 
      x02bai <= 32'b00111111110101010101011110001111;
      x02jyou <= 32'b00111111001100011100101011010010;
    end else if (wbdata[22:12] == 410) begin 
      x02bai <= 32'b00111111110101010100000101011000;
      x02jyou <= 32'b00111111001100011010010111001101;
    end else if (wbdata[22:12] == 411) begin 
      x02bai <= 32'b00111111110101010010101100100101;
      x02jyou <= 32'b00111111001100011000000011010011;
    end else if (wbdata[22:12] == 412) begin 
      x02bai <= 32'b00111111110101010001010011111000;
      x02jyou <= 32'b00111111001100010101101111100110;
    end else if (wbdata[22:12] == 413) begin 
      x02bai <= 32'b00111111110101001111111011001110;
      x02jyou <= 32'b00111111001100010011011100000011;
    end else if (wbdata[22:12] == 414) begin 
      x02bai <= 32'b00111111110101001110100010101010;
      x02jyou <= 32'b00111111001100010001001000101101;
    end else if (wbdata[22:12] == 415) begin 
      x02bai <= 32'b00111111110101001101001010001010;
      x02jyou <= 32'b00111111001100001110110101100010;
    end else if (wbdata[22:12] == 416) begin 
      x02bai <= 32'b00111111110101001011110001101110;
      x02jyou <= 32'b00111111001100001100100010100001;
    end else if (wbdata[22:12] == 417) begin 
      x02bai <= 32'b00111111110101001010011001011000;
      x02jyou <= 32'b00111111001100001010001111101110;
    end else if (wbdata[22:12] == 418) begin 
      x02bai <= 32'b00111111110101001001000001000101;
      x02jyou <= 32'b00111111001100000111111101000100;
    end else if (wbdata[22:12] == 419) begin 
      x02bai <= 32'b00111111110101000111101000111000;
      x02jyou <= 32'b00111111001100000101101010100111;
    end else if (wbdata[22:12] == 420) begin 
      x02bai <= 32'b00111111110101000110010000101111;
      x02jyou <= 32'b00111111001100000011011000010101;
    end else if (wbdata[22:12] == 421) begin 
      x02bai <= 32'b00111111110101000100111000101010;
      x02jyou <= 32'b00111111001100000001000110001101;
    end else if (wbdata[22:12] == 422) begin 
      x02bai <= 32'b00111111110101000011100000101010;
      x02jyou <= 32'b00111111001011111110110100010010;
    end else if (wbdata[22:12] == 423) begin 
      x02bai <= 32'b00111111110101000010001000101111;
      x02jyou <= 32'b00111111001011111100100010100010;
    end else if (wbdata[22:12] == 424) begin 
      x02bai <= 32'b00111111110101000000110000111000;
      x02jyou <= 32'b00111111001011111010010000111101;
    end else if (wbdata[22:12] == 425) begin 
      x02bai <= 32'b00111111110100111111011001000110;
      x02jyou <= 32'b00111111001011110111111111100100;
    end else if (wbdata[22:12] == 426) begin 
      x02bai <= 32'b00111111110100111110000001011000;
      x02jyou <= 32'b00111111001011110101101110010110;
    end else if (wbdata[22:12] == 427) begin 
      x02bai <= 32'b00111111110100111100101001101111;
      x02jyou <= 32'b00111111001011110011011101010011;
    end else if (wbdata[22:12] == 428) begin 
      x02bai <= 32'b00111111110100111011010010001010;
      x02jyou <= 32'b00111111001011110001001100011011;
    end else if (wbdata[22:12] == 429) begin 
      x02bai <= 32'b00111111110100111001111010101010;
      x02jyou <= 32'b00111111001011101110111011101111;
    end else if (wbdata[22:12] == 430) begin 
      x02bai <= 32'b00111111110100111000100011001111;
      x02jyou <= 32'b00111111001011101100101011001110;
    end else if (wbdata[22:12] == 431) begin 
      x02bai <= 32'b00111111110100110111001011111000;
      x02jyou <= 32'b00111111001011101010011010111000;
    end else if (wbdata[22:12] == 432) begin 
      x02bai <= 32'b00111111110100110101110100100101;
      x02jyou <= 32'b00111111001011101000001010101101;
    end else if (wbdata[22:12] == 433) begin 
      x02bai <= 32'b00111111110100110100011101010111;
      x02jyou <= 32'b00111111001011100101111010101101;
    end else if (wbdata[22:12] == 434) begin 
      x02bai <= 32'b00111111110100110011000110001101;
      x02jyou <= 32'b00111111001011100011101010111000;
    end else if (wbdata[22:12] == 435) begin 
      x02bai <= 32'b00111111110100110001101111001000;
      x02jyou <= 32'b00111111001011100001011011001111;
    end else if (wbdata[22:12] == 436) begin 
      x02bai <= 32'b00111111110100110000011000001000;
      x02jyou <= 32'b00111111001011011111001011110001;
    end else if (wbdata[22:12] == 437) begin 
      x02bai <= 32'b00111111110100101111000001001100;
      x02jyou <= 32'b00111111001011011100111100011110;
    end else if (wbdata[22:12] == 438) begin 
      x02bai <= 32'b00111111110100101101101010010100;
      x02jyou <= 32'b00111111001011011010101101010101;
    end else if (wbdata[22:12] == 439) begin 
      x02bai <= 32'b00111111110100101100010011100001;
      x02jyou <= 32'b00111111001011011000011110011001;
    end else if (wbdata[22:12] == 440) begin 
      x02bai <= 32'b00111111110100101010111100110010;
      x02jyou <= 32'b00111111001011010110001111100110;
    end else if (wbdata[22:12] == 441) begin 
      x02bai <= 32'b00111111110100101001100110001000;
      x02jyou <= 32'b00111111001011010100000000111111;
    end else if (wbdata[22:12] == 442) begin 
      x02bai <= 32'b00111111110100101000001111100010;
      x02jyou <= 32'b00111111001011010001110010100011;
    end else if (wbdata[22:12] == 443) begin 
      x02bai <= 32'b00111111110100100110111001000001;
      x02jyou <= 32'b00111111001011001111100100010010;
    end else if (wbdata[22:12] == 444) begin 
      x02bai <= 32'b00111111110100100101100010100100;
      x02jyou <= 32'b00111111001011001101010110001100;
    end else if (wbdata[22:12] == 445) begin 
      x02bai <= 32'b00111111110100100100001100001011;
      x02jyou <= 32'b00111111001011001011001000010000;
    end else if (wbdata[22:12] == 446) begin 
      x02bai <= 32'b00111111110100100010110101110111;
      x02jyou <= 32'b00111111001011001000111010011111;
    end else if (wbdata[22:12] == 447) begin 
      x02bai <= 32'b00111111110100100001011111101000;
      x02jyou <= 32'b00111111001011000110101100111011;
    end else if (wbdata[22:12] == 448) begin 
      x02bai <= 32'b00111111110100100000001001011100;
      x02jyou <= 32'b00111111001011000100011111011111;
    end else if (wbdata[22:12] == 449) begin 
      x02bai <= 32'b00111111110100011110110011010110;
      x02jyou <= 32'b00111111001011000010010010010001;
    end else if (wbdata[22:12] == 450) begin 
      x02bai <= 32'b00111111110100011101011101010011;
      x02jyou <= 32'b00111111001011000000000101001011;
    end else if (wbdata[22:12] == 451) begin 
      x02bai <= 32'b00111111110100011100000111010101;
      x02jyou <= 32'b00111111001010111101111000010001;
    end else if (wbdata[22:12] == 452) begin 
      x02bai <= 32'b00111111110100011010110001011100;
      x02jyou <= 32'b00111111001010111011101011100010;
    end else if (wbdata[22:12] == 453) begin 
      x02bai <= 32'b00111111110100011001011011100111;
      x02jyou <= 32'b00111111001010111001011110111110;
    end else if (wbdata[22:12] == 454) begin 
      x02bai <= 32'b00111111110100011000000101110110;
      x02jyou <= 32'b00111111001010110111010010100100;
    end else if (wbdata[22:12] == 455) begin 
      x02bai <= 32'b00111111110100010110110000001001;
      x02jyou <= 32'b00111111001010110101000110010100;
    end else if (wbdata[22:12] == 456) begin 
      x02bai <= 32'b00111111110100010101011010100001;
      x02jyou <= 32'b00111111001010110010111010010000;
    end else if (wbdata[22:12] == 457) begin 
      x02bai <= 32'b00111111110100010100000100111110;
      x02jyou <= 32'b00111111001010110000101110011000;
    end else if (wbdata[22:12] == 458) begin 
      x02bai <= 32'b00111111110100010010101111011110;
      x02jyou <= 32'b00111111001010101110100010101000;
    end else if (wbdata[22:12] == 459) begin 
      x02bai <= 32'b00111111110100010001011010000100;
      x02jyou <= 32'b00111111001010101100010111000110;
    end else if (wbdata[22:12] == 460) begin 
      x02bai <= 32'b00111111110100010000000100101101;
      x02jyou <= 32'b00111111001010101010001011101011;
    end else if (wbdata[22:12] == 461) begin 
      x02bai <= 32'b00111111110100001110101111011011;
      x02jyou <= 32'b00111111001010101000000000011101;
    end else if (wbdata[22:12] == 462) begin 
      x02bai <= 32'b00111111110100001101011010001101;
      x02jyou <= 32'b00111111001010100101110101011001;
    end else if (wbdata[22:12] == 463) begin 
      x02bai <= 32'b00111111110100001100000101000011;
      x02jyou <= 32'b00111111001010100011101010011111;
    end else if (wbdata[22:12] == 464) begin 
      x02bai <= 32'b00111111110100001010101111111110;
      x02jyou <= 32'b00111111001010100001011111110000;
    end else if (wbdata[22:12] == 465) begin 
      x02bai <= 32'b00111111110100001001011010111101;
      x02jyou <= 32'b00111111001010011111010101001100;
    end else if (wbdata[22:12] == 466) begin 
      x02bai <= 32'b00111111110100001000000110000001;
      x02jyou <= 32'b00111111001010011101001010110011;
    end else if (wbdata[22:12] == 467) begin 
      x02bai <= 32'b00111111110100000110110001001001;
      x02jyou <= 32'b00111111001010011011000000100100;
    end else if (wbdata[22:12] == 468) begin 
      x02bai <= 32'b00111111110100000101011100010101;
      x02jyou <= 32'b00111111001010011000110110100000;
    end else if (wbdata[22:12] == 469) begin 
      x02bai <= 32'b00111111110100000100000111100101;
      x02jyou <= 32'b00111111001010010110101100100101;
    end else if (wbdata[22:12] == 470) begin 
      x02bai <= 32'b00111111110100000010110010111010;
      x02jyou <= 32'b00111111001010010100100010110110;
    end else if (wbdata[22:12] == 471) begin 
      x02bai <= 32'b00111111110100000001011110010011;
      x02jyou <= 32'b00111111001010010010011001010001;
    end else if (wbdata[22:12] == 472) begin 
      x02bai <= 32'b00111111110100000000001001110001;
      x02jyou <= 32'b00111111001010010000001111111000;
    end else if (wbdata[22:12] == 473) begin 
      x02bai <= 32'b00111111110011111110110101010010;
      x02jyou <= 32'b00111111001010001110000110100111;
    end else if (wbdata[22:12] == 474) begin 
      x02bai <= 32'b00111111110011111101100000111000;
      x02jyou <= 32'b00111111001010001011111101100001;
    end else if (wbdata[22:12] == 475) begin 
      x02bai <= 32'b00111111110011111100001100100010;
      x02jyou <= 32'b00111111001010001001110100100110;
    end else if (wbdata[22:12] == 476) begin 
      x02bai <= 32'b00111111110011111010111000010001;
      x02jyou <= 32'b00111111001010000111101011110110;
    end else if (wbdata[22:12] == 477) begin 
      x02bai <= 32'b00111111110011111001100100000100;
      x02jyou <= 32'b00111111001010000101100011010000;
    end else if (wbdata[22:12] == 478) begin 
      x02bai <= 32'b00111111110011111000001111111011;
      x02jyou <= 32'b00111111001010000011011010110100;
    end else if (wbdata[22:12] == 479) begin 
      x02bai <= 32'b00111111110011110110111011110110;
      x02jyou <= 32'b00111111001010000001010010100010;
    end else if (wbdata[22:12] == 480) begin 
      x02bai <= 32'b00111111110011110101100111110101;
      x02jyou <= 32'b00111111001001111111001010011010;
    end else if (wbdata[22:12] == 481) begin 
      x02bai <= 32'b00111111110011110100010011111001;
      x02jyou <= 32'b00111111001001111101000010011101;
    end else if (wbdata[22:12] == 482) begin 
      x02bai <= 32'b00111111110011110011000000000001;
      x02jyou <= 32'b00111111001001111010111010101011;
    end else if (wbdata[22:12] == 483) begin 
      x02bai <= 32'b00111111110011110001101100001110;
      x02jyou <= 32'b00111111001001111000110011000011;
    end else if (wbdata[22:12] == 484) begin 
      x02bai <= 32'b00111111110011110000011000011110;
      x02jyou <= 32'b00111111001001110110101011100101;
    end else if (wbdata[22:12] == 485) begin 
      x02bai <= 32'b00111111110011101111000100110011;
      x02jyou <= 32'b00111111001001110100100100010001;
    end else if (wbdata[22:12] == 486) begin 
      x02bai <= 32'b00111111110011101101110001001100;
      x02jyou <= 32'b00111111001001110010011101001000;
    end else if (wbdata[22:12] == 487) begin 
      x02bai <= 32'b00111111110011101100011101101001;
      x02jyou <= 32'b00111111001001110000010110001000;
    end else if (wbdata[22:12] == 488) begin 
      x02bai <= 32'b00111111110011101011001010001010;
      x02jyou <= 32'b00111111001001101110001111010011;
    end else if (wbdata[22:12] == 489) begin 
      x02bai <= 32'b00111111110011101001110110110000;
      x02jyou <= 32'b00111111001001101100001000101000;
    end else if (wbdata[22:12] == 490) begin 
      x02bai <= 32'b00111111110011101000100011011010;
      x02jyou <= 32'b00111111001001101010000010001000;
    end else if (wbdata[22:12] == 491) begin 
      x02bai <= 32'b00111111110011100111010000001000;
      x02jyou <= 32'b00111111001001100111111011110001;
    end else if (wbdata[22:12] == 492) begin 
      x02bai <= 32'b00111111110011100101111100111010;
      x02jyou <= 32'b00111111001001100101110101100101;
    end else if (wbdata[22:12] == 493) begin 
      x02bai <= 32'b00111111110011100100101001110001;
      x02jyou <= 32'b00111111001001100011101111100100;
    end else if (wbdata[22:12] == 494) begin 
      x02bai <= 32'b00111111110011100011010110101011;
      x02jyou <= 32'b00111111001001100001101001101010;
    end else if (wbdata[22:12] == 495) begin 
      x02bai <= 32'b00111111110011100010000011101010;
      x02jyou <= 32'b00111111001001011111100011111101;
    end else if (wbdata[22:12] == 496) begin 
      x02bai <= 32'b00111111110011100000110000101101;
      x02jyou <= 32'b00111111001001011101011110011001;
    end else if (wbdata[22:12] == 497) begin 
      x02bai <= 32'b00111111110011011111011101110100;
      x02jyou <= 32'b00111111001001011011011000111111;
    end else if (wbdata[22:12] == 498) begin 
      x02bai <= 32'b00111111110011011110001010111111;
      x02jyou <= 32'b00111111001001011001010011101111;
    end else if (wbdata[22:12] == 499) begin 
      x02bai <= 32'b00111111110011011100111000001111;
      x02jyou <= 32'b00111111001001010111001110101010;
    end else if (wbdata[22:12] == 500) begin 
      x02bai <= 32'b00111111110011011011100101100011;
      x02jyou <= 32'b00111111001001010101001001101111;
    end else if (wbdata[22:12] == 501) begin 
      x02bai <= 32'b00111111110011011010010010111010;
      x02jyou <= 32'b00111111001001010011000100111100;
    end else if (wbdata[22:12] == 502) begin 
      x02bai <= 32'b00111111110011011001000000010110;
      x02jyou <= 32'b00111111001001010001000000010100;
    end else if (wbdata[22:12] == 503) begin 
      x02bai <= 32'b00111111110011010111101101110110;
      x02jyou <= 32'b00111111001001001110111011110111;
    end else if (wbdata[22:12] == 504) begin 
      x02bai <= 32'b00111111110011010110011011011010;
      x02jyou <= 32'b00111111001001001100110111100010;
    end else if (wbdata[22:12] == 505) begin 
      x02bai <= 32'b00111111110011010101001001000011;
      x02jyou <= 32'b00111111001001001010110011011010;
    end else if (wbdata[22:12] == 506) begin 
      x02bai <= 32'b00111111110011010011110110101111;
      x02jyou <= 32'b00111111001001001000101111011001;
    end else if (wbdata[22:12] == 507) begin 
      x02bai <= 32'b00111111110011010010100100100000;
      x02jyou <= 32'b00111111001001000110101011100100;
    end else if (wbdata[22:12] == 508) begin 
      x02bai <= 32'b00111111110011010001010010010101;
      x02jyou <= 32'b00111111001001000100100111111000;
    end else if (wbdata[22:12] == 509) begin 
      x02bai <= 32'b00111111110011010000000000001101;
      x02jyou <= 32'b00111111001001000010100100010101;
    end else if (wbdata[22:12] == 510) begin 
      x02bai <= 32'b00111111110011001110101110001010;
      x02jyou <= 32'b00111111001001000000100000111101;
    end else if (wbdata[22:12] == 511) begin 
      x02bai <= 32'b00111111110011001101011100001011;
      x02jyou <= 32'b00111111001000111110011101101110;
    end else if (wbdata[22:12] == 512) begin 
      x02bai <= 32'b00111111110011001100001010010000;
      x02jyou <= 32'b00111111001000111100011010101001;
    end else if (wbdata[22:12] == 513) begin 
      x02bai <= 32'b00111111110011001010111000011010;
      x02jyou <= 32'b00111111001000111010010111110000;
    end else if (wbdata[22:12] == 514) begin 
      x02bai <= 32'b00111111110011001001100110100111;
      x02jyou <= 32'b00111111001000111000010100111110;
    end else if (wbdata[22:12] == 515) begin 
      x02bai <= 32'b00111111110011001000010100111000;
      x02jyou <= 32'b00111111001000110110010010010111;
    end else if (wbdata[22:12] == 516) begin 
      x02bai <= 32'b00111111110011000111000011001110;
      x02jyou <= 32'b00111111001000110100001111111010;
    end else if (wbdata[22:12] == 517) begin 
      x02bai <= 32'b00111111110011000101110001100111;
      x02jyou <= 32'b00111111001000110010001101100110;
    end else if (wbdata[22:12] == 518) begin 
      x02bai <= 32'b00111111110011000100100000000101;
      x02jyou <= 32'b00111111001000110000001011011100;
    end else if (wbdata[22:12] == 519) begin 
      x02bai <= 32'b00111111110011000011001110100111;
      x02jyou <= 32'b00111111001000101110001001011101;
    end else if (wbdata[22:12] == 520) begin 
      x02bai <= 32'b00111111110011000001111101001100;
      x02jyou <= 32'b00111111001000101100000111100101;
    end else if (wbdata[22:12] == 521) begin 
      x02bai <= 32'b00111111110011000000101011110110;
      x02jyou <= 32'b00111111001000101010000101111001;
    end else if (wbdata[22:12] == 522) begin 
      x02bai <= 32'b00111111110010111111011010100100;
      x02jyou <= 32'b00111111001000101000000100010110;
    end else if (wbdata[22:12] == 523) begin 
      x02bai <= 32'b00111111110010111110001001010110;
      x02jyou <= 32'b00111111001000100110000010111100;
    end else if (wbdata[22:12] == 524) begin 
      x02bai <= 32'b00111111110010111100111000001100;
      x02jyou <= 32'b00111111001000100100000001101101;
    end else if (wbdata[22:12] == 525) begin 
      x02bai <= 32'b00111111110010111011100111000110;
      x02jyou <= 32'b00111111001000100010000000100111;
    end else if (wbdata[22:12] == 526) begin 
      x02bai <= 32'b00111111110010111010010110000100;
      x02jyou <= 32'b00111111001000011111111111101010;
    end else if (wbdata[22:12] == 527) begin 
      x02bai <= 32'b00111111110010111001000101000110;
      x02jyou <= 32'b00111111001000011101111110110111;
    end else if (wbdata[22:12] == 528) begin 
      x02bai <= 32'b00111111110010110111110100001100;
      x02jyou <= 32'b00111111001000011011111110001110;
    end else if (wbdata[22:12] == 529) begin 
      x02bai <= 32'b00111111110010110110100011010110;
      x02jyou <= 32'b00111111001000011001111101101110;
    end else if (wbdata[22:12] == 530) begin 
      x02bai <= 32'b00111111110010110101010010100100;
      x02jyou <= 32'b00111111001000010111111101011000;
    end else if (wbdata[22:12] == 531) begin 
      x02bai <= 32'b00111111110010110100000001110110;
      x02jyou <= 32'b00111111001000010101111101001011;
    end else if (wbdata[22:12] == 532) begin 
      x02bai <= 32'b00111111110010110010110001001100;
      x02jyou <= 32'b00111111001000010011111101001000;
    end else if (wbdata[22:12] == 533) begin 
      x02bai <= 32'b00111111110010110001100000100110;
      x02jyou <= 32'b00111111001000010001111101001111;
    end else if (wbdata[22:12] == 534) begin 
      x02bai <= 32'b00111111110010110000010000000100;
      x02jyou <= 32'b00111111001000001111111101011110;
    end else if (wbdata[22:12] == 535) begin 
      x02bai <= 32'b00111111110010101110111111100110;
      x02jyou <= 32'b00111111001000001101111101111000;
    end else if (wbdata[22:12] == 536) begin 
      x02bai <= 32'b00111111110010101101101111001100;
      x02jyou <= 32'b00111111001000001011111110011011;
    end else if (wbdata[22:12] == 537) begin 
      x02bai <= 32'b00111111110010101100011110110110;
      x02jyou <= 32'b00111111001000001001111111000111;
    end else if (wbdata[22:12] == 538) begin 
      x02bai <= 32'b00111111110010101011001110100100;
      x02jyou <= 32'b00111111001000000111111111111101;
    end else if (wbdata[22:12] == 539) begin 
      x02bai <= 32'b00111111110010101001111110010110;
      x02jyou <= 32'b00111111001000000110000000111100;
    end else if (wbdata[22:12] == 540) begin 
      x02bai <= 32'b00111111110010101000101110001100;
      x02jyou <= 32'b00111111001000000100000010000101;
    end else if (wbdata[22:12] == 541) begin 
      x02bai <= 32'b00111111110010100111011110000110;
      x02jyou <= 32'b00111111001000000010000011010111;
    end else if (wbdata[22:12] == 542) begin 
      x02bai <= 32'b00111111110010100110001110000100;
      x02jyou <= 32'b00111111001000000000000100110011;
    end else if (wbdata[22:12] == 543) begin 
      x02bai <= 32'b00111111110010100100111110000110;
      x02jyou <= 32'b00111111000111111110000110011000;
    end else if (wbdata[22:12] == 544) begin 
      x02bai <= 32'b00111111110010100011101110001100;
      x02jyou <= 32'b00111111000111111100001000000111;
    end else if (wbdata[22:12] == 545) begin 
      x02bai <= 32'b00111111110010100010011110010101;
      x02jyou <= 32'b00111111000111111010001001111101;
    end else if (wbdata[22:12] == 546) begin 
      x02bai <= 32'b00111111110010100001001110100011;
      x02jyou <= 32'b00111111000111111000001011111111;
    end else if (wbdata[22:12] == 547) begin 
      x02bai <= 32'b00111111110010011111111110110101;
      x02jyou <= 32'b00111111000111110110001110001010;
    end else if (wbdata[22:12] == 548) begin 
      x02bai <= 32'b00111111110010011110101111001010;
      x02jyou <= 32'b00111111000111110100010000011100;
    end else if (wbdata[22:12] == 549) begin 
      x02bai <= 32'b00111111110010011101011111100100;
      x02jyou <= 32'b00111111000111110010010010111010;
    end else if (wbdata[22:12] == 550) begin 
      x02bai <= 32'b00111111110010011100010000000001;
      x02jyou <= 32'b00111111000111110000010101100000;
    end else if (wbdata[22:12] == 551) begin 
      x02bai <= 32'b00111111110010011011000000100010;
      x02jyou <= 32'b00111111000111101110011000001111;
    end else if (wbdata[22:12] == 552) begin 
      x02bai <= 32'b00111111110010011001110001001000;
      x02jyou <= 32'b00111111000111101100011011001000;
    end else if (wbdata[22:12] == 553) begin 
      x02bai <= 32'b00111111110010011000100001110001;
      x02jyou <= 32'b00111111000111101010011110001010;
    end else if (wbdata[22:12] == 554) begin 
      x02bai <= 32'b00111111110010010111010010011110;
      x02jyou <= 32'b00111111000111101000100001010101;
    end else if (wbdata[22:12] == 555) begin 
      x02bai <= 32'b00111111110010010110000011001111;
      x02jyou <= 32'b00111111000111100110100100101010;
    end else if (wbdata[22:12] == 556) begin 
      x02bai <= 32'b00111111110010010100110100000011;
      x02jyou <= 32'b00111111000111100100101000000110;
    end else if (wbdata[22:12] == 557) begin 
      x02bai <= 32'b00111111110010010011100100111100;
      x02jyou <= 32'b00111111000111100010101011101101;
    end else if (wbdata[22:12] == 558) begin 
      x02bai <= 32'b00111111110010010010010101111001;
      x02jyou <= 32'b00111111000111100000101111011101;
    end else if (wbdata[22:12] == 559) begin 
      x02bai <= 32'b00111111110010010001000110111001;
      x02jyou <= 32'b00111111000111011110110011010110;
    end else if (wbdata[22:12] == 560) begin 
      x02bai <= 32'b00111111110010001111110111111101;
      x02jyou <= 32'b00111111000111011100110111010111;
    end else if (wbdata[22:12] == 561) begin 
      x02bai <= 32'b00111111110010001110101001000110;
      x02jyou <= 32'b00111111000111011010111011100100;
    end else if (wbdata[22:12] == 562) begin 
      x02bai <= 32'b00111111110010001101011010010010;
      x02jyou <= 32'b00111111000111011000111111111000;
    end else if (wbdata[22:12] == 563) begin 
      x02bai <= 32'b00111111110010001100001011100010;
      x02jyou <= 32'b00111111000111010111000100010101;
    end else if (wbdata[22:12] == 564) begin 
      x02bai <= 32'b00111111110010001010111100110101;
      x02jyou <= 32'b00111111000111010101001000111011;
    end else if (wbdata[22:12] == 565) begin 
      x02bai <= 32'b00111111110010001001101110001101;
      x02jyou <= 32'b00111111000111010011001101101011;
    end else if (wbdata[22:12] == 566) begin 
      x02bai <= 32'b00111111110010001000011111101001;
      x02jyou <= 32'b00111111000111010001010010100100;
    end else if (wbdata[22:12] == 567) begin 
      x02bai <= 32'b00111111110010000111010001001000;
      x02jyou <= 32'b00111111000111001111010111100101;
    end else if (wbdata[22:12] == 568) begin 
      x02bai <= 32'b00111111110010000110000010101011;
      x02jyou <= 32'b00111111000111001101011100110000;
    end else if (wbdata[22:12] == 569) begin 
      x02bai <= 32'b00111111110010000100110100010010;
      x02jyou <= 32'b00111111000111001011100010000011;
    end else if (wbdata[22:12] == 570) begin 
      x02bai <= 32'b00111111110010000011100101111101;
      x02jyou <= 32'b00111111000111001001100111100000;
    end else if (wbdata[22:12] == 571) begin 
      x02bai <= 32'b00111111110010000010010111101100;
      x02jyou <= 32'b00111111000111000111101101000110;
    end else if (wbdata[22:12] == 572) begin 
      x02bai <= 32'b00111111110010000001001001011110;
      x02jyou <= 32'b00111111000111000101110010110100;
    end else if (wbdata[22:12] == 573) begin 
      x02bai <= 32'b00111111110001111111111011010100;
      x02jyou <= 32'b00111111000111000011111000101011;
    end else if (wbdata[22:12] == 574) begin 
      x02bai <= 32'b00111111110001111110101101001111;
      x02jyou <= 32'b00111111000111000001111110101101;
    end else if (wbdata[22:12] == 575) begin 
      x02bai <= 32'b00111111110001111101011111001101;
      x02jyou <= 32'b00111111000111000000000100110111;
    end else if (wbdata[22:12] == 576) begin 
      x02bai <= 32'b00111111110001111100010001001110;
      x02jyou <= 32'b00111111000110111110001011001000;
    end else if (wbdata[22:12] == 577) begin 
      x02bai <= 32'b00111111110001111011000011010100;
      x02jyou <= 32'b00111111000110111100010001100100;
    end else if (wbdata[22:12] == 578) begin 
      x02bai <= 32'b00111111110001111001110101011101;
      x02jyou <= 32'b00111111000110111010011000000111;
    end else if (wbdata[22:12] == 579) begin 
      x02bai <= 32'b00111111110001111000100111101010;
      x02jyou <= 32'b00111111000110111000011110110100;
    end else if (wbdata[22:12] == 580) begin 
      x02bai <= 32'b00111111110001110111011001111011;
      x02jyou <= 32'b00111111000110110110100101101010;
    end else if (wbdata[22:12] == 581) begin 
      x02bai <= 32'b00111111110001110110001100010000;
      x02jyou <= 32'b00111111000110110100101100101001;
    end else if (wbdata[22:12] == 582) begin 
      x02bai <= 32'b00111111110001110100111110101000;
      x02jyou <= 32'b00111111000110110010110011110000;
    end else if (wbdata[22:12] == 583) begin 
      x02bai <= 32'b00111111110001110011110001000101;
      x02jyou <= 32'b00111111000110110000111011000001;
    end else if (wbdata[22:12] == 584) begin 
      x02bai <= 32'b00111111110001110010100011100101;
      x02jyou <= 32'b00111111000110101111000010011011;
    end else if (wbdata[22:12] == 585) begin 
      x02bai <= 32'b00111111110001110001010110001001;
      x02jyou <= 32'b00111111000110101101001001111101;
    end else if (wbdata[22:12] == 586) begin 
      x02bai <= 32'b00111111110001110000001000110000;
      x02jyou <= 32'b00111111000110101011010001100111;
    end else if (wbdata[22:12] == 587) begin 
      x02bai <= 32'b00111111110001101110111011011100;
      x02jyou <= 32'b00111111000110101001011001011011;
    end else if (wbdata[22:12] == 588) begin 
      x02bai <= 32'b00111111110001101101101110001011;
      x02jyou <= 32'b00111111000110100111100001010111;
    end else if (wbdata[22:12] == 589) begin 
      x02bai <= 32'b00111111110001101100100000111101;
      x02jyou <= 32'b00111111000110100101101001011011;
    end else if (wbdata[22:12] == 590) begin 
      x02bai <= 32'b00111111110001101011010011110100;
      x02jyou <= 32'b00111111000110100011110001101001;
    end else if (wbdata[22:12] == 591) begin 
      x02bai <= 32'b00111111110001101010000110101110;
      x02jyou <= 32'b00111111000110100001111001111111;
    end else if (wbdata[22:12] == 592) begin 
      x02bai <= 32'b00111111110001101000111001101100;
      x02jyou <= 32'b00111111000110100000000010011110;
    end else if (wbdata[22:12] == 593) begin 
      x02bai <= 32'b00111111110001100111101100101110;
      x02jyou <= 32'b00111111000110011110001011000110;
    end else if (wbdata[22:12] == 594) begin 
      x02bai <= 32'b00111111110001100110011111110100;
      x02jyou <= 32'b00111111000110011100010011111000;
    end else if (wbdata[22:12] == 595) begin 
      x02bai <= 32'b00111111110001100101010010111101;
      x02jyou <= 32'b00111111000110011010011100110000;
    end else if (wbdata[22:12] == 596) begin 
      x02bai <= 32'b00111111110001100100000110001010;
      x02jyou <= 32'b00111111000110011000100101110010;
    end else if (wbdata[22:12] == 597) begin 
      x02bai <= 32'b00111111110001100010111001011011;
      x02jyou <= 32'b00111111000110010110101110111101;
    end else if (wbdata[22:12] == 598) begin 
      x02bai <= 32'b00111111110001100001101100101111;
      x02jyou <= 32'b00111111000110010100111000010000;
    end else if (wbdata[22:12] == 599) begin 
      x02bai <= 32'b00111111110001100000100000000111;
      x02jyou <= 32'b00111111000110010011000001101011;
    end else if (wbdata[22:12] == 600) begin 
      x02bai <= 32'b00111111110001011111010011100011;
      x02jyou <= 32'b00111111000110010001001011010000;
    end else if (wbdata[22:12] == 601) begin 
      x02bai <= 32'b00111111110001011110000111000010;
      x02jyou <= 32'b00111111000110001111010100111100;
    end else if (wbdata[22:12] == 602) begin 
      x02bai <= 32'b00111111110001011100111010100110;
      x02jyou <= 32'b00111111000110001101011110110010;
    end else if (wbdata[22:12] == 603) begin 
      x02bai <= 32'b00111111110001011011101110001100;
      x02jyou <= 32'b00111111000110001011101000101111;
    end else if (wbdata[22:12] == 604) begin 
      x02bai <= 32'b00111111110001011010100001110111;
      x02jyou <= 32'b00111111000110001001110010110110;
    end else if (wbdata[22:12] == 605) begin 
      x02bai <= 32'b00111111110001011001010101100101;
      x02jyou <= 32'b00111111000110000111111101000101;
    end else if (wbdata[22:12] == 606) begin 
      x02bai <= 32'b00111111110001011000001001010111;
      x02jyou <= 32'b00111111000110000110000111011100;
    end else if (wbdata[22:12] == 607) begin 
      x02bai <= 32'b00111111110001010110111101001101;
      x02jyou <= 32'b00111111000110000100010001111101;
    end else if (wbdata[22:12] == 608) begin 
      x02bai <= 32'b00111111110001010101110001000110;
      x02jyou <= 32'b00111111000110000010011100100101;
    end else if (wbdata[22:12] == 609) begin 
      x02bai <= 32'b00111111110001010100100101000011;
      x02jyou <= 32'b00111111000110000000100111010110;
    end else if (wbdata[22:12] == 610) begin 
      x02bai <= 32'b00111111110001010011011001000100;
      x02jyou <= 32'b00111111000101111110110010010000;
    end else if (wbdata[22:12] == 611) begin 
      x02bai <= 32'b00111111110001010010001101001000;
      x02jyou <= 32'b00111111000101111100111101010010;
    end else if (wbdata[22:12] == 612) begin 
      x02bai <= 32'b00111111110001010001000001010000;
      x02jyou <= 32'b00111111000101111011001000011100;
    end else if (wbdata[22:12] == 613) begin 
      x02bai <= 32'b00111111110001001111110101011011;
      x02jyou <= 32'b00111111000101111001010011101110;
    end else if (wbdata[22:12] == 614) begin 
      x02bai <= 32'b00111111110001001110101001101011;
      x02jyou <= 32'b00111111000101110111011111001010;
    end else if (wbdata[22:12] == 615) begin 
      x02bai <= 32'b00111111110001001101011101111101;
      x02jyou <= 32'b00111111000101110101101010101101;
    end else if (wbdata[22:12] == 616) begin 
      x02bai <= 32'b00111111110001001100010010010100;
      x02jyou <= 32'b00111111000101110011110110011010;
    end else if (wbdata[22:12] == 617) begin 
      x02bai <= 32'b00111111110001001011000110101110;
      x02jyou <= 32'b00111111000101110010000010001110;
    end else if (wbdata[22:12] == 618) begin 
      x02bai <= 32'b00111111110001001001111011001100;
      x02jyou <= 32'b00111111000101110000001110001011;
    end else if (wbdata[22:12] == 619) begin 
      x02bai <= 32'b00111111110001001000101111101101;
      x02jyou <= 32'b00111111000101101110011010001111;
    end else if (wbdata[22:12] == 620) begin 
      x02bai <= 32'b00111111110001000111100100010010;
      x02jyou <= 32'b00111111000101101100100110011101;
    end else if (wbdata[22:12] == 621) begin 
      x02bai <= 32'b00111111110001000110011000111011;
      x02jyou <= 32'b00111111000101101010110010110011;
    end else if (wbdata[22:12] == 622) begin 
      x02bai <= 32'b00111111110001000101001101100111;
      x02jyou <= 32'b00111111000101101000111111010001;
    end else if (wbdata[22:12] == 623) begin 
      x02bai <= 32'b00111111110001000100000010010111;
      x02jyou <= 32'b00111111000101100111001011111000;
    end else if (wbdata[22:12] == 624) begin 
      x02bai <= 32'b00111111110001000010110111001010;
      x02jyou <= 32'b00111111000101100101011000100110;
    end else if (wbdata[22:12] == 625) begin 
      x02bai <= 32'b00111111110001000001101100000001;
      x02jyou <= 32'b00111111000101100011100101011100;
    end else if (wbdata[22:12] == 626) begin 
      x02bai <= 32'b00111111110001000000100000111100;
      x02jyou <= 32'b00111111000101100001110010011100;
    end else if (wbdata[22:12] == 627) begin 
      x02bai <= 32'b00111111110000111111010101111010;
      x02jyou <= 32'b00111111000101011111111111100011;
    end else if (wbdata[22:12] == 628) begin 
      x02bai <= 32'b00111111110000111110001010111100;
      x02jyou <= 32'b00111111000101011110001100110011;
    end else if (wbdata[22:12] == 629) begin 
      x02bai <= 32'b00111111110000111101000000000001;
      x02jyou <= 32'b00111111000101011100011010001011;
    end else if (wbdata[22:12] == 630) begin 
      x02bai <= 32'b00111111110000111011110101001010;
      x02jyou <= 32'b00111111000101011010100111101011;
    end else if (wbdata[22:12] == 631) begin 
      x02bai <= 32'b00111111110000111010101010010111;
      x02jyou <= 32'b00111111000101011000110101010100;
    end else if (wbdata[22:12] == 632) begin 
      x02bai <= 32'b00111111110000111001011111100111;
      x02jyou <= 32'b00111111000101010111000011000100;
    end else if (wbdata[22:12] == 633) begin 
      x02bai <= 32'b00111111110000111000010100111011;
      x02jyou <= 32'b00111111000101010101010000111101;
    end else if (wbdata[22:12] == 634) begin 
      x02bai <= 32'b00111111110000110111001010010010;
      x02jyou <= 32'b00111111000101010011011110111110;
    end else if (wbdata[22:12] == 635) begin 
      x02bai <= 32'b00111111110000110101111111101101;
      x02jyou <= 32'b00111111000101010001101101000111;
    end else if (wbdata[22:12] == 636) begin 
      x02bai <= 32'b00111111110000110100110101001011;
      x02jyou <= 32'b00111111000101001111111011011000;
    end else if (wbdata[22:12] == 637) begin 
      x02bai <= 32'b00111111110000110011101010101101;
      x02jyou <= 32'b00111111000101001110001001110001;
    end else if (wbdata[22:12] == 638) begin 
      x02bai <= 32'b00111111110000110010100000010010;
      x02jyou <= 32'b00111111000101001100011000010010;
    end else if (wbdata[22:12] == 639) begin 
      x02bai <= 32'b00111111110000110001010101111011;
      x02jyou <= 32'b00111111000101001010100110111011;
    end else if (wbdata[22:12] == 640) begin 
      x02bai <= 32'b00111111110000110000001011101000;
      x02jyou <= 32'b00111111000101001000110101101101;
    end else if (wbdata[22:12] == 641) begin 
      x02bai <= 32'b00111111110000101111000001011000;
      x02jyou <= 32'b00111111000101000111000100100111;
    end else if (wbdata[22:12] == 642) begin 
      x02bai <= 32'b00111111110000101101110111001100;
      x02jyou <= 32'b00111111000101000101010011101001;
    end else if (wbdata[22:12] == 643) begin 
      x02bai <= 32'b00111111110000101100101101000011;
      x02jyou <= 32'b00111111000101000011100010110011;
    end else if (wbdata[22:12] == 644) begin 
      x02bai <= 32'b00111111110000101011100010111101;
      x02jyou <= 32'b00111111000101000001110010000100;
    end else if (wbdata[22:12] == 645) begin 
      x02bai <= 32'b00111111110000101010011000111100;
      x02jyou <= 32'b00111111000101000000000001011111;
    end else if (wbdata[22:12] == 646) begin 
      x02bai <= 32'b00111111110000101001001110111101;
      x02jyou <= 32'b00111111000100111110010001000000;
    end else if (wbdata[22:12] == 647) begin 
      x02bai <= 32'b00111111110000101000000101000011;
      x02jyou <= 32'b00111111000100111100100000101011;
    end else if (wbdata[22:12] == 648) begin 
      x02bai <= 32'b00111111110000100110111011001011;
      x02jyou <= 32'b00111111000100111010110000011100;
    end else if (wbdata[22:12] == 649) begin 
      x02bai <= 32'b00111111110000100101110001011000;
      x02jyou <= 32'b00111111000100111001000000010111;
    end else if (wbdata[22:12] == 650) begin 
      x02bai <= 32'b00111111110000100100100111100111;
      x02jyou <= 32'b00111111000100110111010000010111;
    end else if (wbdata[22:12] == 651) begin 
      x02bai <= 32'b00111111110000100011011101111011;
      x02jyou <= 32'b00111111000100110101100000100010;
    end else if (wbdata[22:12] == 652) begin 
      x02bai <= 32'b00111111110000100010010100010001;
      x02jyou <= 32'b00111111000100110011110000110011;
    end else if (wbdata[22:12] == 653) begin 
      x02bai <= 32'b00111111110000100001001010101011;
      x02jyou <= 32'b00111111000100110010000001001101;
    end else if (wbdata[22:12] == 654) begin 
      x02bai <= 32'b00111111110000100000000001001001;
      x02jyou <= 32'b00111111000100110000010001101111;
    end else if (wbdata[22:12] == 655) begin 
      x02bai <= 32'b00111111110000011110110111101010;
      x02jyou <= 32'b00111111000100101110100010011000;
    end else if (wbdata[22:12] == 656) begin 
      x02bai <= 32'b00111111110000011101101110001111;
      x02jyou <= 32'b00111111000100101100110011001010;
    end else if (wbdata[22:12] == 657) begin 
      x02bai <= 32'b00111111110000011100100100110111;
      x02jyou <= 32'b00111111000100101011000100000011;
    end else if (wbdata[22:12] == 658) begin 
      x02bai <= 32'b00111111110000011011011011100011;
      x02jyou <= 32'b00111111000100101001010101000101;
    end else if (wbdata[22:12] == 659) begin 
      x02bai <= 32'b00111111110000011010010010010010;
      x02jyou <= 32'b00111111000100100111100110001110;
    end else if (wbdata[22:12] == 660) begin 
      x02bai <= 32'b00111111110000011001001001000100;
      x02jyou <= 32'b00111111000100100101110111011110;
    end else if (wbdata[22:12] == 661) begin 
      x02bai <= 32'b00111111110000010111111111111010;
      x02jyou <= 32'b00111111000100100100001000110111;
    end else if (wbdata[22:12] == 662) begin 
      x02bai <= 32'b00111111110000010110110110110100;
      x02jyou <= 32'b00111111000100100010011010011000;
    end else if (wbdata[22:12] == 663) begin 
      x02bai <= 32'b00111111110000010101101101110001;
      x02jyou <= 32'b00111111000100100000101100000001;
    end else if (wbdata[22:12] == 664) begin 
      x02bai <= 32'b00111111110000010100100100110001;
      x02jyou <= 32'b00111111000100011110111101110001;
    end else if (wbdata[22:12] == 665) begin 
      x02bai <= 32'b00111111110000010011011011110101;
      x02jyou <= 32'b00111111000100011101001111101001;
    end else if (wbdata[22:12] == 666) begin 
      x02bai <= 32'b00111111110000010010010010111100;
      x02jyou <= 32'b00111111000100011011100001101001;
    end else if (wbdata[22:12] == 667) begin 
      x02bai <= 32'b00111111110000010001001010000111;
      x02jyou <= 32'b00111111000100011001110011110001;
    end else if (wbdata[22:12] == 668) begin 
      x02bai <= 32'b00111111110000010000000001010101;
      x02jyou <= 32'b00111111000100011000000110000000;
    end else if (wbdata[22:12] == 669) begin 
      x02bai <= 32'b00111111110000001110111000100110;
      x02jyou <= 32'b00111111000100010110011000010111;
    end else if (wbdata[22:12] == 670) begin 
      x02bai <= 32'b00111111110000001101101111111011;
      x02jyou <= 32'b00111111000100010100101010110110;
    end else if (wbdata[22:12] == 671) begin 
      x02bai <= 32'b00111111110000001100100111010100;
      x02jyou <= 32'b00111111000100010010111101011101;
    end else if (wbdata[22:12] == 672) begin 
      x02bai <= 32'b00111111110000001011011110110000;
      x02jyou <= 32'b00111111000100010001010000001100;
    end else if (wbdata[22:12] == 673) begin 
      x02bai <= 32'b00111111110000001010010110001111;
      x02jyou <= 32'b00111111000100001111100011000010;
    end else if (wbdata[22:12] == 674) begin 
      x02bai <= 32'b00111111110000001001001101110001;
      x02jyou <= 32'b00111111000100001101110101111110;
    end else if (wbdata[22:12] == 675) begin 
      x02bai <= 32'b00111111110000001000000101010111;
      x02jyou <= 32'b00111111000100001100001001000100;
    end else if (wbdata[22:12] == 676) begin 
      x02bai <= 32'b00111111110000000110111101000001;
      x02jyou <= 32'b00111111000100001010011100010010;
    end else if (wbdata[22:12] == 677) begin 
      x02bai <= 32'b00111111110000000101110100101110;
      x02jyou <= 32'b00111111000100001000101111100111;
    end else if (wbdata[22:12] == 678) begin 
      x02bai <= 32'b00111111110000000100101100011110;
      x02jyou <= 32'b00111111000100000111000011000011;
    end else if (wbdata[22:12] == 679) begin 
      x02bai <= 32'b00111111110000000011100100010001;
      x02jyou <= 32'b00111111000100000101010110100110;
    end else if (wbdata[22:12] == 680) begin 
      x02bai <= 32'b00111111110000000010011100001000;
      x02jyou <= 32'b00111111000100000011101010010010;
    end else if (wbdata[22:12] == 681) begin 
      x02bai <= 32'b00111111110000000001010100000011;
      x02jyou <= 32'b00111111000100000001111110000110;
    end else if (wbdata[22:12] == 682) begin 
      x02bai <= 32'b00111111110000000000001100000000;
      x02jyou <= 32'b00111111000100000000010010000000;
    end else if (wbdata[22:12] == 683) begin 
      x02bai <= 32'b00111111101111111111000100000010;
      x02jyou <= 32'b00111111000011111110100110000100;
    end else if (wbdata[22:12] == 684) begin 
      x02bai <= 32'b00111111101111111101111100000110;
      x02jyou <= 32'b00111111000011111100111010001101;
    end else if (wbdata[22:12] == 685) begin 
      x02bai <= 32'b00111111101111111100110100001110;
      x02jyou <= 32'b00111111000011111011001110011111;
    end else if (wbdata[22:12] == 686) begin 
      x02bai <= 32'b00111111101111111011101100011001;
      x02jyou <= 32'b00111111000011111001100010111000;
    end else if (wbdata[22:12] == 687) begin 
      x02bai <= 32'b00111111101111111010100100101000;
      x02jyou <= 32'b00111111000011110111110111011001;
    end else if (wbdata[22:12] == 688) begin 
      x02bai <= 32'b00111111101111111001011100111010;
      x02jyou <= 32'b00111111000011110110001100000010;
    end else if (wbdata[22:12] == 689) begin 
      x02bai <= 32'b00111111101111111000010101001111;
      x02jyou <= 32'b00111111000011110100100000110001;
    end else if (wbdata[22:12] == 690) begin 
      x02bai <= 32'b00111111101111110111001101101000;
      x02jyou <= 32'b00111111000011110010110101101001;
    end else if (wbdata[22:12] == 691) begin 
      x02bai <= 32'b00111111101111110110000110000100;
      x02jyou <= 32'b00111111000011110001001010101000;
    end else if (wbdata[22:12] == 692) begin 
      x02bai <= 32'b00111111101111110100111110100011;
      x02jyou <= 32'b00111111000011101111011111101110;
    end else if (wbdata[22:12] == 693) begin 
      x02bai <= 32'b00111111101111110011110111000110;
      x02jyou <= 32'b00111111000011101101110100111100;
    end else if (wbdata[22:12] == 694) begin 
      x02bai <= 32'b00111111101111110010101111101100;
      x02jyou <= 32'b00111111000011101100001010010010;
    end else if (wbdata[22:12] == 695) begin 
      x02bai <= 32'b00111111101111110001101000010101;
      x02jyou <= 32'b00111111000011101010011111101110;
    end else if (wbdata[22:12] == 696) begin 
      x02bai <= 32'b00111111101111110000100001000010;
      x02jyou <= 32'b00111111000011101000110101010011;
    end else if (wbdata[22:12] == 697) begin 
      x02bai <= 32'b00111111101111101111011001110010;
      x02jyou <= 32'b00111111000011100111001010111110;
    end else if (wbdata[22:12] == 698) begin 
      x02bai <= 32'b00111111101111101110010010100101;
      x02jyou <= 32'b00111111000011100101100000110001;
    end else if (wbdata[22:12] == 699) begin 
      x02bai <= 32'b00111111101111101101001011011100;
      x02jyou <= 32'b00111111000011100011110110101100;
    end else if (wbdata[22:12] == 700) begin 
      x02bai <= 32'b00111111101111101100000100010110;
      x02jyou <= 32'b00111111000011100010001100101110;
    end else if (wbdata[22:12] == 701) begin 
      x02bai <= 32'b00111111101111101010111101010011;
      x02jyou <= 32'b00111111000011100000100010110111;
    end else if (wbdata[22:12] == 702) begin 
      x02bai <= 32'b00111111101111101001110110010011;
      x02jyou <= 32'b00111111000011011110111001000111;
    end else if (wbdata[22:12] == 703) begin 
      x02bai <= 32'b00111111101111101000101111010111;
      x02jyou <= 32'b00111111000011011101001111100000;
    end else if (wbdata[22:12] == 704) begin 
      x02bai <= 32'b00111111101111100111101000011110;
      x02jyou <= 32'b00111111000011011011100101111111;
    end else if (wbdata[22:12] == 705) begin 
      x02bai <= 32'b00111111101111100110100001101001;
      x02jyou <= 32'b00111111000011011001111100100110;
    end else if (wbdata[22:12] == 706) begin 
      x02bai <= 32'b00111111101111100101011010110111;
      x02jyou <= 32'b00111111000011011000010011010101;
    end else if (wbdata[22:12] == 707) begin 
      x02bai <= 32'b00111111101111100100010100001000;
      x02jyou <= 32'b00111111000011010110101010001010;
    end else if (wbdata[22:12] == 708) begin 
      x02bai <= 32'b00111111101111100011001101011100;
      x02jyou <= 32'b00111111000011010101000001000111;
    end else if (wbdata[22:12] == 709) begin 
      x02bai <= 32'b00111111101111100010000110110100;
      x02jyou <= 32'b00111111000011010011011000001100;
    end else if (wbdata[22:12] == 710) begin 
      x02bai <= 32'b00111111101111100001000000001111;
      x02jyou <= 32'b00111111000011010001101111010111;
    end else if (wbdata[22:12] == 711) begin 
      x02bai <= 32'b00111111101111011111111001101101;
      x02jyou <= 32'b00111111000011010000000110101010;
    end else if (wbdata[22:12] == 712) begin 
      x02bai <= 32'b00111111101111011110110011001110;
      x02jyou <= 32'b00111111000011001110011110000011;
    end else if (wbdata[22:12] == 713) begin 
      x02bai <= 32'b00111111101111011101101100110011;
      x02jyou <= 32'b00111111000011001100110101100101;
    end else if (wbdata[22:12] == 714) begin 
      x02bai <= 32'b00111111101111011100100110011011;
      x02jyou <= 32'b00111111000011001011001101001110;
    end else if (wbdata[22:12] == 715) begin 
      x02bai <= 32'b00111111101111011011100000000110;
      x02jyou <= 32'b00111111000011001001100100111101;
    end else if (wbdata[22:12] == 716) begin 
      x02bai <= 32'b00111111101111011010011001110100;
      x02jyou <= 32'b00111111000011000111111100110100;
    end else if (wbdata[22:12] == 717) begin 
      x02bai <= 32'b00111111101111011001010011100110;
      x02jyou <= 32'b00111111000011000110010100110010;
    end else if (wbdata[22:12] == 718) begin 
      x02bai <= 32'b00111111101111011000001101011011;
      x02jyou <= 32'b00111111000011000100101100111000;
    end else if (wbdata[22:12] == 719) begin 
      x02bai <= 32'b00111111101111010111000111010011;
      x02jyou <= 32'b00111111000011000011000101000100;
    end else if (wbdata[22:12] == 720) begin 
      x02bai <= 32'b00111111101111010110000001001111;
      x02jyou <= 32'b00111111000011000001011101011001;
    end else if (wbdata[22:12] == 721) begin 
      x02bai <= 32'b00111111101111010100111011001110;
      x02jyou <= 32'b00111111000010111111110101110100;
    end else if (wbdata[22:12] == 722) begin 
      x02bai <= 32'b00111111101111010011110101001111;
      x02jyou <= 32'b00111111000010111110001110010101;
    end else if (wbdata[22:12] == 723) begin 
      x02bai <= 32'b00111111101111010010101111010101;
      x02jyou <= 32'b00111111000010111100100111000000;
    end else if (wbdata[22:12] == 724) begin 
      x02bai <= 32'b00111111101111010001101001011101;
      x02jyou <= 32'b00111111000010111010111111110000;
    end else if (wbdata[22:12] == 725) begin 
      x02bai <= 32'b00111111101111010000100011101001;
      x02jyou <= 32'b00111111000010111001011000101000;
    end else if (wbdata[22:12] == 726) begin 
      x02bai <= 32'b00111111101111001111011101110111;
      x02jyou <= 32'b00111111000010110111110001100110;
    end else if (wbdata[22:12] == 727) begin 
      x02bai <= 32'b00111111101111001110011000001010;
      x02jyou <= 32'b00111111000010110110001010101101;
    end else if (wbdata[22:12] == 728) begin 
      x02bai <= 32'b00111111101111001101010010011111;
      x02jyou <= 32'b00111111000010110100100011111010;
    end else if (wbdata[22:12] == 729) begin 
      x02bai <= 32'b00111111101111001100001100110111;
      x02jyou <= 32'b00111111000010110010111101001110;
    end else if (wbdata[22:12] == 730) begin 
      x02bai <= 32'b00111111101111001011000111010011;
      x02jyou <= 32'b00111111000010110001010110101001;
    end else if (wbdata[22:12] == 731) begin 
      x02bai <= 32'b00111111101111001010000001110010;
      x02jyou <= 32'b00111111000010101111110000001100;
    end else if (wbdata[22:12] == 732) begin 
      x02bai <= 32'b00111111101111001000111100010100;
      x02jyou <= 32'b00111111000010101110001001110101;
    end else if (wbdata[22:12] == 733) begin 
      x02bai <= 32'b00111111101111000111110110111001;
      x02jyou <= 32'b00111111000010101100100011100101;
    end else if (wbdata[22:12] == 734) begin 
      x02bai <= 32'b00111111101111000110110001100010;
      x02jyou <= 32'b00111111000010101010111101011110;
    end else if (wbdata[22:12] == 735) begin 
      x02bai <= 32'b00111111101111000101101100001101;
      x02jyou <= 32'b00111111000010101001010111011011;
    end else if (wbdata[22:12] == 736) begin 
      x02bai <= 32'b00111111101111000100100110111100;
      x02jyou <= 32'b00111111000010100111110001100001;
    end else if (wbdata[22:12] == 737) begin 
      x02bai <= 32'b00111111101111000011100001101110;
      x02jyou <= 32'b00111111000010100110001011101110;
    end else if (wbdata[22:12] == 738) begin 
      x02bai <= 32'b00111111101111000010011100100100;
      x02jyou <= 32'b00111111000010100100100110000011;
    end else if (wbdata[22:12] == 739) begin 
      x02bai <= 32'b00111111101111000001010111011100;
      x02jyou <= 32'b00111111000010100011000000011101;
    end else if (wbdata[22:12] == 740) begin 
      x02bai <= 32'b00111111101111000000010010011000;
      x02jyou <= 32'b00111111000010100001011010111111;
    end else if (wbdata[22:12] == 741) begin 
      x02bai <= 32'b00111111101110111111001101010110;
      x02jyou <= 32'b00111111000010011111110101100111;
    end else if (wbdata[22:12] == 742) begin 
      x02bai <= 32'b00111111101110111110001000011000;
      x02jyou <= 32'b00111111000010011110010000010111;
    end else if (wbdata[22:12] == 743) begin 
      x02bai <= 32'b00111111101110111101000011011101;
      x02jyou <= 32'b00111111000010011100101011001101;
    end else if (wbdata[22:12] == 744) begin 
      x02bai <= 32'b00111111101110111011111110100101;
      x02jyou <= 32'b00111111000010011011000110001011;
    end else if (wbdata[22:12] == 745) begin 
      x02bai <= 32'b00111111101110111010111001110001;
      x02jyou <= 32'b00111111000010011001100001010000;
    end else if (wbdata[22:12] == 746) begin 
      x02bai <= 32'b00111111101110111001110100111111;
      x02jyou <= 32'b00111111000010010111111100011011;
    end else if (wbdata[22:12] == 747) begin 
      x02bai <= 32'b00111111101110111000110000010001;
      x02jyou <= 32'b00111111000010010110010111101101;
    end else if (wbdata[22:12] == 748) begin 
      x02bai <= 32'b00111111101110110111101011100110;
      x02jyou <= 32'b00111111000010010100110011000111;
    end else if (wbdata[22:12] == 749) begin 
      x02bai <= 32'b00111111101110110110100110111110;
      x02jyou <= 32'b00111111000010010011001110100111;
    end else if (wbdata[22:12] == 750) begin 
      x02bai <= 32'b00111111101110110101100010011001;
      x02jyou <= 32'b00111111000010010001101010001110;
    end else if (wbdata[22:12] == 751) begin 
      x02bai <= 32'b00111111101110110100011101110111;
      x02jyou <= 32'b00111111000010010000000101111100;
    end else if (wbdata[22:12] == 752) begin 
      x02bai <= 32'b00111111101110110011011001011001;
      x02jyou <= 32'b00111111000010001110100001110010;
    end else if (wbdata[22:12] == 753) begin 
      x02bai <= 32'b00111111101110110010010100111101;
      x02jyou <= 32'b00111111000010001100111101101101;
    end else if (wbdata[22:12] == 754) begin 
      x02bai <= 32'b00111111101110110001010000100101;
      x02jyou <= 32'b00111111000010001011011001110000;
    end else if (wbdata[22:12] == 755) begin 
      x02bai <= 32'b00111111101110110000001100010000;
      x02jyou <= 32'b00111111000010001001110101111001;
    end else if (wbdata[22:12] == 756) begin 
      x02bai <= 32'b00111111101110101111000111111101;
      x02jyou <= 32'b00111111000010001000010010001000;
    end else if (wbdata[22:12] == 757) begin 
      x02bai <= 32'b00111111101110101110000011101110;
      x02jyou <= 32'b00111111000010000110101110011111;
    end else if (wbdata[22:12] == 758) begin 
      x02bai <= 32'b00111111101110101100111111100010;
      x02jyou <= 32'b00111111000010000101001010111101;
    end else if (wbdata[22:12] == 759) begin 
      x02bai <= 32'b00111111101110101011111011011010;
      x02jyou <= 32'b00111111000010000011100111100011;
    end else if (wbdata[22:12] == 760) begin 
      x02bai <= 32'b00111111101110101010110111010100;
      x02jyou <= 32'b00111111000010000010000100001110;
    end else if (wbdata[22:12] == 761) begin 
      x02bai <= 32'b00111111101110101001110011010001;
      x02jyou <= 32'b00111111000010000000100001000000;
    end else if (wbdata[22:12] == 762) begin 
      x02bai <= 32'b00111111101110101000101111010010;
      x02jyou <= 32'b00111111000001111110111101111010;
    end else if (wbdata[22:12] == 763) begin 
      x02bai <= 32'b00111111101110100111101011010110;
      x02jyou <= 32'b00111111000001111101011010111010;
    end else if (wbdata[22:12] == 764) begin 
      x02bai <= 32'b00111111101110100110100111011100;
      x02jyou <= 32'b00111111000001111011110111111111;
    end else if (wbdata[22:12] == 765) begin 
      x02bai <= 32'b00111111101110100101100011100110;
      x02jyou <= 32'b00111111000001111010010101001101;
    end else if (wbdata[22:12] == 766) begin 
      x02bai <= 32'b00111111101110100100011111110011;
      x02jyou <= 32'b00111111000001111000110010100001;
    end else if (wbdata[22:12] == 767) begin 
      x02bai <= 32'b00111111101110100011011100000011;
      x02jyou <= 32'b00111111000001110111001111111100;
    end else if (wbdata[22:12] == 768) begin 
      x02bai <= 32'b00111111101110100010011000010110;
      x02jyou <= 32'b00111111000001110101101101011110;
    end else if (wbdata[22:12] == 769) begin 
      x02bai <= 32'b00111111101110100001010100101100;
      x02jyou <= 32'b00111111000001110100001011000110;
    end else if (wbdata[22:12] == 770) begin 
      x02bai <= 32'b00111111101110100000010001000101;
      x02jyou <= 32'b00111111000001110010101000110100;
    end else if (wbdata[22:12] == 771) begin 
      x02bai <= 32'b00111111101110011111001101100001;
      x02jyou <= 32'b00111111000001110001000110101010;
    end else if (wbdata[22:12] == 772) begin 
      x02bai <= 32'b00111111101110011110001010000001;
      x02jyou <= 32'b00111111000001101111100100100111;
    end else if (wbdata[22:12] == 773) begin 
      x02bai <= 32'b00111111101110011101000110100011;
      x02jyou <= 32'b00111111000001101110000010101001;
    end else if (wbdata[22:12] == 774) begin 
      x02bai <= 32'b00111111101110011100000011001001;
      x02jyou <= 32'b00111111000001101100100000110100;
    end else if (wbdata[22:12] == 775) begin 
      x02bai <= 32'b00111111101110011010111111110001;
      x02jyou <= 32'b00111111000001101010111111000011;
    end else if (wbdata[22:12] == 776) begin 
      x02bai <= 32'b00111111101110011001111100011101;
      x02jyou <= 32'b00111111000001101001011101011011;
    end else if (wbdata[22:12] == 777) begin 
      x02bai <= 32'b00111111101110011000111001001011;
      x02jyou <= 32'b00111111000001100111111011110111;
    end else if (wbdata[22:12] == 778) begin 
      x02bai <= 32'b00111111101110010111110101111101;
      x02jyou <= 32'b00111111000001100110011010011100;
    end else if (wbdata[22:12] == 779) begin 
      x02bai <= 32'b00111111101110010110110010110010;
      x02jyou <= 32'b00111111000001100100111001000111;
    end else if (wbdata[22:12] == 780) begin 
      x02bai <= 32'b00111111101110010101101111101001;
      x02jyou <= 32'b00111111000001100011010111111000;
    end else if (wbdata[22:12] == 781) begin 
      x02bai <= 32'b00111111101110010100101100100100;
      x02jyou <= 32'b00111111000001100001110110110000;
    end else if (wbdata[22:12] == 782) begin 
      x02bai <= 32'b00111111101110010011101001100010;
      x02jyou <= 32'b00111111000001100000010101101111;
    end else if (wbdata[22:12] == 783) begin 
      x02bai <= 32'b00111111101110010010100110100011;
      x02jyou <= 32'b00111111000001011110110100110100;
    end else if (wbdata[22:12] == 784) begin 
      x02bai <= 32'b00111111101110010001100011100111;
      x02jyou <= 32'b00111111000001011101010100000000;
    end else if (wbdata[22:12] == 785) begin 
      x02bai <= 32'b00111111101110010000100000101110;
      x02jyou <= 32'b00111111000001011011110011010011;
    end else if (wbdata[22:12] == 786) begin 
      x02bai <= 32'b00111111101110001111011101110111;
      x02jyou <= 32'b00111111000001011010010010101010;
    end else if (wbdata[22:12] == 787) begin 
      x02bai <= 32'b00111111101110001110011011000100;
      x02jyou <= 32'b00111111000001011000110010001010;
    end else if (wbdata[22:12] == 788) begin 
      x02bai <= 32'b00111111101110001101011000010100;
      x02jyou <= 32'b00111111000001010111010001110000;
    end else if (wbdata[22:12] == 789) begin 
      x02bai <= 32'b00111111101110001100010101100111;
      x02jyou <= 32'b00111111000001010101110001011100;
    end else if (wbdata[22:12] == 790) begin 
      x02bai <= 32'b00111111101110001011010010111101;
      x02jyou <= 32'b00111111000001010100010001001111;
    end else if (wbdata[22:12] == 791) begin 
      x02bai <= 32'b00111111101110001010010000010110;
      x02jyou <= 32'b00111111000001010010110001001001;
    end else if (wbdata[22:12] == 792) begin 
      x02bai <= 32'b00111111101110001001001101110010;
      x02jyou <= 32'b00111111000001010001010001001001;
    end else if (wbdata[22:12] == 793) begin 
      x02bai <= 32'b00111111101110001000001011010001;
      x02jyou <= 32'b00111111000001001111110001001111;
    end else if (wbdata[22:12] == 794) begin 
      x02bai <= 32'b00111111101110000111001000110011;
      x02jyou <= 32'b00111111000001001110010001011100;
    end else if (wbdata[22:12] == 795) begin 
      x02bai <= 32'b00111111101110000110000110011000;
      x02jyou <= 32'b00111111000001001100110001110000;
    end else if (wbdata[22:12] == 796) begin 
      x02bai <= 32'b00111111101110000101000100000000;
      x02jyou <= 32'b00111111000001001011010010001010;
    end else if (wbdata[22:12] == 797) begin 
      x02bai <= 32'b00111111101110000100000001101011;
      x02jyou <= 32'b00111111000001001001110010101010;
    end else if (wbdata[22:12] == 798) begin 
      x02bai <= 32'b00111111101110000010111111011001;
      x02jyou <= 32'b00111111000001001000010011010001;
    end else if (wbdata[22:12] == 799) begin 
      x02bai <= 32'b00111111101110000001111101001010;
      x02jyou <= 32'b00111111000001000110110011111110;
    end else if (wbdata[22:12] == 800) begin 
      x02bai <= 32'b00111111101110000000111010111110;
      x02jyou <= 32'b00111111000001000101010100110010;
    end else if (wbdata[22:12] == 801) begin 
      x02bai <= 32'b00111111101101111111111000110100;
      x02jyou <= 32'b00111111000001000011110101101011;
    end else if (wbdata[22:12] == 802) begin 
      x02bai <= 32'b00111111101101111110110110101110;
      x02jyou <= 32'b00111111000001000010010110101011;
    end else if (wbdata[22:12] == 803) begin 
      x02bai <= 32'b00111111101101111101110100101011;
      x02jyou <= 32'b00111111000001000000110111110011;
    end else if (wbdata[22:12] == 804) begin 
      x02bai <= 32'b00111111101101111100110010101011;
      x02jyou <= 32'b00111111000000111111011001000000;
    end else if (wbdata[22:12] == 805) begin 
      x02bai <= 32'b00111111101101111011110000101101;
      x02jyou <= 32'b00111111000000111101111010010011;
    end else if (wbdata[22:12] == 806) begin 
      x02bai <= 32'b00111111101101111010101110110011;
      x02jyou <= 32'b00111111000000111100011011101101;
    end else if (wbdata[22:12] == 807) begin 
      x02bai <= 32'b00111111101101111001101100111100;
      x02jyou <= 32'b00111111000000111010111101001110;
    end else if (wbdata[22:12] == 808) begin 
      x02bai <= 32'b00111111101101111000101011000111;
      x02jyou <= 32'b00111111000000111001011110110100;
    end else if (wbdata[22:12] == 809) begin 
      x02bai <= 32'b00111111101101110111101001010110;
      x02jyou <= 32'b00111111000000111000000000100001;
    end else if (wbdata[22:12] == 810) begin 
      x02bai <= 32'b00111111101101110110100111100111;
      x02jyou <= 32'b00111111000000110110100010010100;
    end else if (wbdata[22:12] == 811) begin 
      x02bai <= 32'b00111111101101110101100101111100;
      x02jyou <= 32'b00111111000000110101000100001111;
    end else if (wbdata[22:12] == 812) begin 
      x02bai <= 32'b00111111101101110100100100010011;
      x02jyou <= 32'b00111111000000110011100110001110;
    end else if (wbdata[22:12] == 813) begin 
      x02bai <= 32'b00111111101101110011100010101101;
      x02jyou <= 32'b00111111000000110010001000010100;
    end else if (wbdata[22:12] == 814) begin 
      x02bai <= 32'b00111111101101110010100001001010;
      x02jyou <= 32'b00111111000000110000101010100000;
    end else if (wbdata[22:12] == 815) begin 
      x02bai <= 32'b00111111101101110001011111101011;
      x02jyou <= 32'b00111111000000101111001100110100;
    end else if (wbdata[22:12] == 816) begin 
      x02bai <= 32'b00111111101101110000011110001110;
      x02jyou <= 32'b00111111000000101101101111001101;
    end else if (wbdata[22:12] == 817) begin 
      x02bai <= 32'b00111111101101101111011100110100;
      x02jyou <= 32'b00111111000000101100010001101101;
    end else if (wbdata[22:12] == 818) begin 
      x02bai <= 32'b00111111101101101110011011011101;
      x02jyou <= 32'b00111111000000101010110100010010;
    end else if (wbdata[22:12] == 819) begin 
      x02bai <= 32'b00111111101101101101011010001000;
      x02jyou <= 32'b00111111000000101001010110111101;
    end else if (wbdata[22:12] == 820) begin 
      x02bai <= 32'b00111111101101101100011000110111;
      x02jyou <= 32'b00111111000000100111111001110000;
    end else if (wbdata[22:12] == 821) begin 
      x02bai <= 32'b00111111101101101011010111101001;
      x02jyou <= 32'b00111111000000100110011100101001;
    end else if (wbdata[22:12] == 822) begin 
      x02bai <= 32'b00111111101101101010010110011101;
      x02jyou <= 32'b00111111000000100100111111100110;
    end else if (wbdata[22:12] == 823) begin 
      x02bai <= 32'b00111111101101101001010101010101;
      x02jyou <= 32'b00111111000000100011100010101100;
    end else if (wbdata[22:12] == 824) begin 
      x02bai <= 32'b00111111101101101000010100001111;
      x02jyou <= 32'b00111111000000100010000101110110;
    end else if (wbdata[22:12] == 825) begin 
      x02bai <= 32'b00111111101101100111010011001100;
      x02jyou <= 32'b00111111000000100000101001000111;
    end else if (wbdata[22:12] == 826) begin 
      x02bai <= 32'b00111111101101100110010010001101;
      x02jyou <= 32'b00111111000000011111001100100000;
    end else if (wbdata[22:12] == 827) begin 
      x02bai <= 32'b00111111101101100101010001010000;
      x02jyou <= 32'b00111111000000011101101111111110;
    end else if (wbdata[22:12] == 828) begin 
      x02bai <= 32'b00111111101101100100010000010110;
      x02jyou <= 32'b00111111000000011100010011100001;
    end else if (wbdata[22:12] == 829) begin 
      x02bai <= 32'b00111111101101100011001111011110;
      x02jyou <= 32'b00111111000000011010110111001010;
    end else if (wbdata[22:12] == 830) begin 
      x02bai <= 32'b00111111101101100010001110101010;
      x02jyou <= 32'b00111111000000011001011010111011;
    end else if (wbdata[22:12] == 831) begin 
      x02bai <= 32'b00111111101101100001001101111001;
      x02jyou <= 32'b00111111000000010111111110110010;
    end else if (wbdata[22:12] == 832) begin 
      x02bai <= 32'b00111111101101100000001101001010;
      x02jyou <= 32'b00111111000000010110100010101101;
    end else if (wbdata[22:12] == 833) begin 
      x02bai <= 32'b00111111101101011111001100011111;
      x02jyou <= 32'b00111111000000010101000110110001;
    end else if (wbdata[22:12] == 834) begin 
      x02bai <= 32'b00111111101101011110001011110110;
      x02jyou <= 32'b00111111000000010011101010111001;
    end else if (wbdata[22:12] == 835) begin 
      x02bai <= 32'b00111111101101011101001011010000;
      x02jyou <= 32'b00111111000000010010001111001000;
    end else if (wbdata[22:12] == 836) begin 
      x02bai <= 32'b00111111101101011100001010101101;
      x02jyou <= 32'b00111111000000010000110011011101;
    end else if (wbdata[22:12] == 837) begin 
      x02bai <= 32'b00111111101101011011001010001101;
      x02jyou <= 32'b00111111000000001111010111111000;
    end else if (wbdata[22:12] == 838) begin 
      x02bai <= 32'b00111111101101011010001001101111;
      x02jyou <= 32'b00111111000000001101111100011000;
    end else if (wbdata[22:12] == 839) begin 
      x02bai <= 32'b00111111101101011001001001010101;
      x02jyou <= 32'b00111111000000001100100001000000;
    end else if (wbdata[22:12] == 840) begin 
      x02bai <= 32'b00111111101101011000001000111101;
      x02jyou <= 32'b00111111000000001011000101101101;
    end else if (wbdata[22:12] == 841) begin 
      x02bai <= 32'b00111111101101010111001000101000;
      x02jyou <= 32'b00111111000000001001101010011111;
    end else if (wbdata[22:12] == 842) begin 
      x02bai <= 32'b00111111101101010110001000010111;
      x02jyou <= 32'b00111111000000001000001111011010;
    end else if (wbdata[22:12] == 843) begin 
      x02bai <= 32'b00111111101101010101001000001000;
      x02jyou <= 32'b00111111000000000110110100011010;
    end else if (wbdata[22:12] == 844) begin 
      x02bai <= 32'b00111111101101010100000111111011;
      x02jyou <= 32'b00111111000000000101011001011110;
    end else if (wbdata[22:12] == 845) begin 
      x02bai <= 32'b00111111101101010011000111110010;
      x02jyou <= 32'b00111111000000000011111110101010;
    end else if (wbdata[22:12] == 846) begin 
      x02bai <= 32'b00111111101101010010000111101011;
      x02jyou <= 32'b00111111000000000010100011111011;
    end else if (wbdata[22:12] == 847) begin 
      x02bai <= 32'b00111111101101010001000111101000;
      x02jyou <= 32'b00111111000000000001001001010011;
    end else if (wbdata[22:12] == 848) begin 
      x02bai <= 32'b00111111101101010000000111100111;
      x02jyou <= 32'b00111110111111111111011101100001;
    end else if (wbdata[22:12] == 849) begin 
      x02bai <= 32'b00111111101101001111000111101001;
      x02jyou <= 32'b00111110111111111100101000101001;
    end else if (wbdata[22:12] == 850) begin 
      x02bai <= 32'b00111111101101001110000111101110;
      x02jyou <= 32'b00111110111111111001110011111100;
    end else if (wbdata[22:12] == 851) begin 
      x02bai <= 32'b00111111101101001101000111110101;
      x02jyou <= 32'b00111110111111110110111111011001;
    end else if (wbdata[22:12] == 852) begin 
      x02bai <= 32'b00111111101101001100001000000000;
      x02jyou <= 32'b00111110111111110100001011000110;
    end else if (wbdata[22:12] == 853) begin 
      x02bai <= 32'b00111111101101001011001000001101;
      x02jyou <= 32'b00111110111111110001010110111100;
    end else if (wbdata[22:12] == 854) begin 
      x02bai <= 32'b00111111101101001010001000011101;
      x02jyou <= 32'b00111110111111101110100010111111;
    end else if (wbdata[22:12] == 855) begin 
      x02bai <= 32'b00111111101101001001001000110000;
      x02jyou <= 32'b00111110111111101011101111001110;
    end else if (wbdata[22:12] == 856) begin 
      x02bai <= 32'b00111111101101001000001001000101;
      x02jyou <= 32'b00111110111111101000111011100111;
    end else if (wbdata[22:12] == 857) begin 
      x02bai <= 32'b00111111101101000111001001011110;
      x02jyou <= 32'b00111110111111100110001000001111;
    end else if (wbdata[22:12] == 858) begin 
      x02bai <= 32'b00111111101101000110001001111001;
      x02jyou <= 32'b00111110111111100011010101000000;
    end else if (wbdata[22:12] == 859) begin 
      x02bai <= 32'b00111111101101000101001010010111;
      x02jyou <= 32'b00111110111111100000100001111110;
    end else if (wbdata[22:12] == 860) begin 
      x02bai <= 32'b00111111101101000100001010111000;
      x02jyou <= 32'b00111110111111011101101111001000;
    end else if (wbdata[22:12] == 861) begin 
      x02bai <= 32'b00111111101101000011001011011100;
      x02jyou <= 32'b00111110111111011010111100011111;
    end else if (wbdata[22:12] == 862) begin 
      x02bai <= 32'b00111111101101000010001100000010;
      x02jyou <= 32'b00111110111111011000001001111111;
    end else if (wbdata[22:12] == 863) begin 
      x02bai <= 32'b00111111101101000001001100101011;
      x02jyou <= 32'b00111110111111010101010111101100;
    end else if (wbdata[22:12] == 864) begin 
      x02bai <= 32'b00111111101101000000001101010111;
      x02jyou <= 32'b00111110111111010010100101100101;
    end else if (wbdata[22:12] == 865) begin 
      x02bai <= 32'b00111111101100111111001110000110;
      x02jyou <= 32'b00111110111111001111110011101010;
    end else if (wbdata[22:12] == 866) begin 
      x02bai <= 32'b00111111101100111110001110111000;
      x02jyou <= 32'b00111110111111001101000001111100;
    end else if (wbdata[22:12] == 867) begin 
      x02bai <= 32'b00111111101100111101001111101100;
      x02jyou <= 32'b00111110111111001010010000010111;
    end else if (wbdata[22:12] == 868) begin 
      x02bai <= 32'b00111111101100111100010000100011;
      x02jyou <= 32'b00111110111111000111011110111110;
    end else if (wbdata[22:12] == 869) begin 
      x02bai <= 32'b00111111101100111011010001011101;
      x02jyou <= 32'b00111110111111000100101101110010;
    end else if (wbdata[22:12] == 870) begin 
      x02bai <= 32'b00111111101100111010010010011010;
      x02jyou <= 32'b00111110111111000001111100110010;
    end else if (wbdata[22:12] == 871) begin 
      x02bai <= 32'b00111111101100111001010011011001;
      x02jyou <= 32'b00111110111110111111001011111100;
    end else if (wbdata[22:12] == 872) begin 
      x02bai <= 32'b00111111101100111000010100011011;
      x02jyou <= 32'b00111110111110111100011011010010;
    end else if (wbdata[22:12] == 873) begin 
      x02bai <= 32'b00111111101100110111010101100000;
      x02jyou <= 32'b00111110111110111001101010110100;
    end else if (wbdata[22:12] == 874) begin 
      x02bai <= 32'b00111111101100110110010110101000;
      x02jyou <= 32'b00111110111110110110111010100011;
    end else if (wbdata[22:12] == 875) begin 
      x02bai <= 32'b00111111101100110101010111110011;
      x02jyou <= 32'b00111110111110110100001010011101;
    end else if (wbdata[22:12] == 876) begin 
      x02bai <= 32'b00111111101100110100011001000000;
      x02jyou <= 32'b00111110111110110001011010100010;
    end else if (wbdata[22:12] == 877) begin 
      x02bai <= 32'b00111111101100110011011010010000;
      x02jyou <= 32'b00111110111110101110101010110010;
    end else if (wbdata[22:12] == 878) begin 
      x02bai <= 32'b00111111101100110010011011100010;
      x02jyou <= 32'b00111110111110101011111011001100;
    end else if (wbdata[22:12] == 879) begin 
      x02bai <= 32'b00111111101100110001011100111000;
      x02jyou <= 32'b00111110111110101001001011110101;
    end else if (wbdata[22:12] == 880) begin 
      x02bai <= 32'b00111111101100110000011110010000;
      x02jyou <= 32'b00111110111110100110011100100111;
    end else if (wbdata[22:12] == 881) begin 
      x02bai <= 32'b00111111101100101111011111101011;
      x02jyou <= 32'b00111110111110100011101101100110;
    end else if (wbdata[22:12] == 882) begin 
      x02bai <= 32'b00111111101100101110100001001001;
      x02jyou <= 32'b00111110111110100000111110110001;
    end else if (wbdata[22:12] == 883) begin 
      x02bai <= 32'b00111111101100101101100010101001;
      x02jyou <= 32'b00111110111110011110010000000101;
    end else if (wbdata[22:12] == 884) begin 
      x02bai <= 32'b00111111101100101100100100001100;
      x02jyou <= 32'b00111110111110011011100001100101;
    end else if (wbdata[22:12] == 885) begin 
      x02bai <= 32'b00111111101100101011100101110010;
      x02jyou <= 32'b00111110111110011000110011010010;
    end else if (wbdata[22:12] == 886) begin 
      x02bai <= 32'b00111111101100101010100111011011;
      x02jyou <= 32'b00111110111110010110000101001010;
    end else if (wbdata[22:12] == 887) begin 
      x02bai <= 32'b00111111101100101001101001000110;
      x02jyou <= 32'b00111110111110010011010111001101;
    end else if (wbdata[22:12] == 888) begin 
      x02bai <= 32'b00111111101100101000101010110100;
      x02jyou <= 32'b00111110111110010000101001011011;
    end else if (wbdata[22:12] == 889) begin 
      x02bai <= 32'b00111111101100100111101100100101;
      x02jyou <= 32'b00111110111110001101111011110101;
    end else if (wbdata[22:12] == 890) begin 
      x02bai <= 32'b00111111101100100110101110011000;
      x02jyou <= 32'b00111110111110001011001110011001;
    end else if (wbdata[22:12] == 891) begin 
      x02bai <= 32'b00111111101100100101110000001110;
      x02jyou <= 32'b00111110111110001000100001001001;
    end else if (wbdata[22:12] == 892) begin 
      x02bai <= 32'b00111111101100100100110010000111;
      x02jyou <= 32'b00111110111110000101110100000101;
    end else if (wbdata[22:12] == 893) begin 
      x02bai <= 32'b00111111101100100011110100000010;
      x02jyou <= 32'b00111110111110000011000111001011;
    end else if (wbdata[22:12] == 894) begin 
      x02bai <= 32'b00111111101100100010110110000001;
      x02jyou <= 32'b00111110111110000000011010011111;
    end else if (wbdata[22:12] == 895) begin 
      x02bai <= 32'b00111111101100100001111000000010;
      x02jyou <= 32'b00111110111101111101101101111101;
    end else if (wbdata[22:12] == 896) begin 
      x02bai <= 32'b00111111101100100000111010000101;
      x02jyou <= 32'b00111110111101111011000001100100;
    end else if (wbdata[22:12] == 897) begin 
      x02bai <= 32'b00111111101100011111111100001100;
      x02jyou <= 32'b00111110111101111000010101011001;
    end else if (wbdata[22:12] == 898) begin 
      x02bai <= 32'b00111111101100011110111110010101;
      x02jyou <= 32'b00111110111101110101101001011001;
    end else if (wbdata[22:12] == 899) begin 
      x02bai <= 32'b00111111101100011110000000100000;
      x02jyou <= 32'b00111110111101110010111101100001;
    end else if (wbdata[22:12] == 900) begin 
      x02bai <= 32'b00111111101100011101000010101111;
      x02jyou <= 32'b00111110111101110000010001111000;
    end else if (wbdata[22:12] == 901) begin 
      x02bai <= 32'b00111111101100011100000101000000;
      x02jyou <= 32'b00111110111101101101100110011001;
    end else if (wbdata[22:12] == 902) begin 
      x02bai <= 32'b00111111101100011011000111010011;
      x02jyou <= 32'b00111110111101101010111011000011;
    end else if (wbdata[22:12] == 903) begin 
      x02bai <= 32'b00111111101100011010001001101010;
      x02jyou <= 32'b00111110111101101000001111111011;
    end else if (wbdata[22:12] == 904) begin 
      x02bai <= 32'b00111111101100011001001100000011;
      x02jyou <= 32'b00111110111101100101100100111101;
    end else if (wbdata[22:12] == 905) begin 
      x02bai <= 32'b00111111101100011000001110011111;
      x02jyou <= 32'b00111110111101100010111010001011;
    end else if (wbdata[22:12] == 906) begin 
      x02bai <= 32'b00111111101100010111010000111101;
      x02jyou <= 32'b00111110111101100000001111100010;
    end else if (wbdata[22:12] == 907) begin 
      x02bai <= 32'b00111111101100010110010011011110;
      x02jyou <= 32'b00111110111101011101100101000101;
    end else if (wbdata[22:12] == 908) begin 
      x02bai <= 32'b00111111101100010101010110000010;
      x02jyou <= 32'b00111110111101011010111010110101;
    end else if (wbdata[22:12] == 909) begin 
      x02bai <= 32'b00111111101100010100011000101000;
      x02jyou <= 32'b00111110111101011000010000101101;
    end else if (wbdata[22:12] == 910) begin 
      x02bai <= 32'b00111111101100010011011011010001;
      x02jyou <= 32'b00111110111101010101100110110001;
    end else if (wbdata[22:12] == 911) begin 
      x02bai <= 32'b00111111101100010010011101111101;
      x02jyou <= 32'b00111110111101010010111101000010;
    end else if (wbdata[22:12] == 912) begin 
      x02bai <= 32'b00111111101100010001100000101100;
      x02jyou <= 32'b00111110111101010000010011011110;
    end else if (wbdata[22:12] == 913) begin 
      x02bai <= 32'b00111111101100010000100011011101;
      x02jyou <= 32'b00111110111101001101101010000100;
    end else if (wbdata[22:12] == 914) begin 
      x02bai <= 32'b00111111101100001111100110010000;
      x02jyou <= 32'b00111110111101001011000000110011;
    end else if (wbdata[22:12] == 915) begin 
      x02bai <= 32'b00111111101100001110101001000111;
      x02jyou <= 32'b00111110111101001000010111110000;
    end else if (wbdata[22:12] == 916) begin 
      x02bai <= 32'b00111111101100001101101100000000;
      x02jyou <= 32'b00111110111101000101101110110111;
    end else if (wbdata[22:12] == 917) begin 
      x02bai <= 32'b00111111101100001100101110111011;
      x02jyou <= 32'b00111110111101000011000110000111;
    end else if (wbdata[22:12] == 918) begin 
      x02bai <= 32'b00111111101100001011110001111001;
      x02jyou <= 32'b00111110111101000000011101100010;
    end else if (wbdata[22:12] == 919) begin 
      x02bai <= 32'b00111111101100001010110100111010;
      x02jyou <= 32'b00111110111100111101110101001010;
    end else if (wbdata[22:12] == 920) begin 
      x02bai <= 32'b00111111101100001001110111111110;
      x02jyou <= 32'b00111110111100111011001100111110;
    end else if (wbdata[22:12] == 921) begin 
      x02bai <= 32'b00111111101100001000111011000100;
      x02jyou <= 32'b00111110111100111000100100111010;
    end else if (wbdata[22:12] == 922) begin 
      x02bai <= 32'b00111111101100000111111110001101;
      x02jyou <= 32'b00111110111100110101111101000011;
    end else if (wbdata[22:12] == 923) begin 
      x02bai <= 32'b00111111101100000111000001011000;
      x02jyou <= 32'b00111110111100110011010101010101;
    end else if (wbdata[22:12] == 924) begin 
      x02bai <= 32'b00111111101100000110000100100110;
      x02jyou <= 32'b00111110111100110000101101110010;
    end else if (wbdata[22:12] == 925) begin 
      x02bai <= 32'b00111111101100000101000111110110;
      x02jyou <= 32'b00111110111100101110000110011001;
    end else if (wbdata[22:12] == 926) begin 
      x02bai <= 32'b00111111101100000100001011001010;
      x02jyou <= 32'b00111110111100101011011111001110;
    end else if (wbdata[22:12] == 927) begin 
      x02bai <= 32'b00111111101100000011001110011111;
      x02jyou <= 32'b00111110111100101000111000001010;
    end else if (wbdata[22:12] == 928) begin 
      x02bai <= 32'b00111111101100000010010001111000;
      x02jyou <= 32'b00111110111100100110010001010100;
    end else if (wbdata[22:12] == 929) begin 
      x02bai <= 32'b00111111101100000001010101010011;
      x02jyou <= 32'b00111110111100100011101010101000;
    end else if (wbdata[22:12] == 930) begin 
      x02bai <= 32'b00111111101100000000011000110001;
      x02jyou <= 32'b00111110111100100001000100000111;
    end else if (wbdata[22:12] == 931) begin 
      x02bai <= 32'b00111111101011111111011100010001;
      x02jyou <= 32'b00111110111100011110011101101111;
    end else if (wbdata[22:12] == 932) begin 
      x02bai <= 32'b00111111101011111110011111110100;
      x02jyou <= 32'b00111110111100011011110111100100;
    end else if (wbdata[22:12] == 933) begin 
      x02bai <= 32'b00111111101011111101100011011001;
      x02jyou <= 32'b00111110111100011001010001100001;
    end else if (wbdata[22:12] == 934) begin 
      x02bai <= 32'b00111111101011111100100111000001;
      x02jyou <= 32'b00111110111100010110101011101010;
    end else if (wbdata[22:12] == 935) begin 
      x02bai <= 32'b00111111101011111011101010101100;
      x02jyou <= 32'b00111110111100010100000101111111;
    end else if (wbdata[22:12] == 936) begin 
      x02bai <= 32'b00111111101011111010101110011001;
      x02jyou <= 32'b00111110111100010001100000011100;
    end else if (wbdata[22:12] == 937) begin 
      x02bai <= 32'b00111111101011111001110010001001;
      x02jyou <= 32'b00111110111100001110111011000110;
    end else if (wbdata[22:12] == 938) begin 
      x02bai <= 32'b00111111101011111000110101111011;
      x02jyou <= 32'b00111110111100001100010101111001;
    end else if (wbdata[22:12] == 939) begin 
      x02bai <= 32'b00111111101011110111111001110000;
      x02jyou <= 32'b00111110111100001001110000110111;
    end else if (wbdata[22:12] == 940) begin 
      x02bai <= 32'b00111111101011110110111101101000;
      x02jyou <= 32'b00111110111100000111001100000001;
    end else if (wbdata[22:12] == 941) begin 
      x02bai <= 32'b00111111101011110110000001100010;
      x02jyou <= 32'b00111110111100000100100111010101;
    end else if (wbdata[22:12] == 942) begin 
      x02bai <= 32'b00111111101011110101000101011110;
      x02jyou <= 32'b00111110111100000010000010110001;
    end else if (wbdata[22:12] == 943) begin 
      x02bai <= 32'b00111111101011110100001001011110;
      x02jyou <= 32'b00111110111011111111011110011011;
    end else if (wbdata[22:12] == 944) begin 
      x02bai <= 32'b00111111101011110011001101011111;
      x02jyou <= 32'b00111110111011111100111010001100;
    end else if (wbdata[22:12] == 945) begin 
      x02bai <= 32'b00111111101011110010010001100100;
      x02jyou <= 32'b00111110111011111010010110001100;
    end else if (wbdata[22:12] == 946) begin 
      x02bai <= 32'b00111111101011110001010101101011;
      x02jyou <= 32'b00111110111011110111110010010100;
    end else if (wbdata[22:12] == 947) begin 
      x02bai <= 32'b00111111101011110000011001110100;
      x02jyou <= 32'b00111110111011110101001110100110;
    end else if (wbdata[22:12] == 948) begin 
      x02bai <= 32'b00111111101011101111011110000000;
      x02jyou <= 32'b00111110111011110010101011000011;
    end else if (wbdata[22:12] == 949) begin 
      x02bai <= 32'b00111111101011101110100010001111;
      x02jyou <= 32'b00111110111011110000000111101011;
    end else if (wbdata[22:12] == 950) begin 
      x02bai <= 32'b00111111101011101101100110100000;
      x02jyou <= 32'b00111110111011101101100100011101;
    end else if (wbdata[22:12] == 951) begin 
      x02bai <= 32'b00111111101011101100101010110100;
      x02jyou <= 32'b00111110111011101011000001011010;
    end else if (wbdata[22:12] == 952) begin 
      x02bai <= 32'b00111111101011101011101111001010;
      x02jyou <= 32'b00111110111011101000011110100001;
    end else if (wbdata[22:12] == 953) begin 
      x02bai <= 32'b00111111101011101010110011100011;
      x02jyou <= 32'b00111110111011100101111011110011;
    end else if (wbdata[22:12] == 954) begin 
      x02bai <= 32'b00111111101011101001110111111110;
      x02jyou <= 32'b00111110111011100011011001001110;
    end else if (wbdata[22:12] == 955) begin 
      x02bai <= 32'b00111111101011101000111100011100;
      x02jyou <= 32'b00111110111011100000110110110100;
    end else if (wbdata[22:12] == 956) begin 
      x02bai <= 32'b00111111101011101000000000111100;
      x02jyou <= 32'b00111110111011011110010100100100;
    end else if (wbdata[22:12] == 957) begin 
      x02bai <= 32'b00111111101011100111000101011111;
      x02jyou <= 32'b00111110111011011011110010011111;
    end else if (wbdata[22:12] == 958) begin 
      x02bai <= 32'b00111111101011100110001010000101;
      x02jyou <= 32'b00111110111011011001010000100101;
    end else if (wbdata[22:12] == 959) begin 
      x02bai <= 32'b00111111101011100101001110101101;
      x02jyou <= 32'b00111110111011010110101110110101;
    end else if (wbdata[22:12] == 960) begin 
      x02bai <= 32'b00111111101011100100010011010111;
      x02jyou <= 32'b00111110111011010100001101001110;
    end else if (wbdata[22:12] == 961) begin 
      x02bai <= 32'b00111111101011100011011000000100;
      x02jyou <= 32'b00111110111011010001101011110010;
    end else if (wbdata[22:12] == 962) begin 
      x02bai <= 32'b00111111101011100010011100110100;
      x02jyou <= 32'b00111110111011001111001010100001;
    end else if (wbdata[22:12] == 963) begin 
      x02bai <= 32'b00111111101011100001100001100110;
      x02jyou <= 32'b00111110111011001100101001011010;
    end else if (wbdata[22:12] == 964) begin 
      x02bai <= 32'b00111111101011100000100110011011;
      x02jyou <= 32'b00111110111011001010001000011110;
    end else if (wbdata[22:12] == 965) begin 
      x02bai <= 32'b00111111101011011111101011010010;
      x02jyou <= 32'b00111110111011000111100111101011;
    end else if (wbdata[22:12] == 966) begin 
      x02bai <= 32'b00111111101011011110110000001011;
      x02jyou <= 32'b00111110111011000101000111000001;
    end else if (wbdata[22:12] == 967) begin 
      x02bai <= 32'b00111111101011011101110101000111;
      x02jyou <= 32'b00111110111011000010100110100010;
    end else if (wbdata[22:12] == 968) begin 
      x02bai <= 32'b00111111101011011100111010000110;
      x02jyou <= 32'b00111110111011000000000110001111;
    end else if (wbdata[22:12] == 969) begin 
      x02bai <= 32'b00111111101011011011111111000111;
      x02jyou <= 32'b00111110111010111101100110000101;
    end else if (wbdata[22:12] == 970) begin 
      x02bai <= 32'b00111111101011011011000100001011;
      x02jyou <= 32'b00111110111010111011000110000111;
    end else if (wbdata[22:12] == 971) begin 
      x02bai <= 32'b00111111101011011010001001010001;
      x02jyou <= 32'b00111110111010111000100110010001;
    end else if (wbdata[22:12] == 972) begin 
      x02bai <= 32'b00111111101011011001001110011010;
      x02jyou <= 32'b00111110111010110110000110100110;
    end else if (wbdata[22:12] == 973) begin 
      x02bai <= 32'b00111111101011011000010011100101;
      x02jyou <= 32'b00111110111010110011100111000101;
    end else if (wbdata[22:12] == 974) begin 
      x02bai <= 32'b00111111101011010111011000110011;
      x02jyou <= 32'b00111110111010110001000111101111;
    end else if (wbdata[22:12] == 975) begin 
      x02bai <= 32'b00111111101011010110011110000011;
      x02jyou <= 32'b00111110111010101110101000100010;
    end else if (wbdata[22:12] == 976) begin 
      x02bai <= 32'b00111111101011010101100011010101;
      x02jyou <= 32'b00111110111010101100001001011101;
    end else if (wbdata[22:12] == 977) begin 
      x02bai <= 32'b00111111101011010100101000101010;
      x02jyou <= 32'b00111110111010101001101010100101;
    end else if (wbdata[22:12] == 978) begin 
      x02bai <= 32'b00111111101011010011101110000010;
      x02jyou <= 32'b00111110111010100111001011110111;
    end else if (wbdata[22:12] == 979) begin 
      x02bai <= 32'b00111111101011010010110011011100;
      x02jyou <= 32'b00111110111010100100101101010010;
    end else if (wbdata[22:12] == 980) begin 
      x02bai <= 32'b00111111101011010001111000111001;
      x02jyou <= 32'b00111110111010100010001110111001;
    end else if (wbdata[22:12] == 981) begin 
      x02bai <= 32'b00111111101011010000111110011000;
      x02jyou <= 32'b00111110111010011111110000101001;
    end else if (wbdata[22:12] == 982) begin 
      x02bai <= 32'b00111111101011010000000011111001;
      x02jyou <= 32'b00111110111010011101010010100001;
    end else if (wbdata[22:12] == 983) begin 
      x02bai <= 32'b00111111101011001111001001011101;
      x02jyou <= 32'b00111110111010011010110100100101;
    end else if (wbdata[22:12] == 984) begin 
      x02bai <= 32'b00111111101011001110001111000011;
      x02jyou <= 32'b00111110111010011000010110110001;
    end else if (wbdata[22:12] == 985) begin 
      x02bai <= 32'b00111111101011001101010100101100;
      x02jyou <= 32'b00111110111010010101111001001001;
    end else if (wbdata[22:12] == 986) begin 
      x02bai <= 32'b00111111101011001100011010011000;
      x02jyou <= 32'b00111110111010010011011011101101;
    end else if (wbdata[22:12] == 987) begin 
      x02bai <= 32'b00111111101011001011100000000101;
      x02jyou <= 32'b00111110111010010000111110010110;
    end else if (wbdata[22:12] == 988) begin 
      x02bai <= 32'b00111111101011001010100101110110;
      x02jyou <= 32'b00111110111010001110100001001101;
    end else if (wbdata[22:12] == 989) begin 
      x02bai <= 32'b00111111101011001001101011101000;
      x02jyou <= 32'b00111110111010001100000100001011;
    end else if (wbdata[22:12] == 990) begin 
      x02bai <= 32'b00111111101011001000110001011101;
      x02jyou <= 32'b00111110111010001001100111010100;
    end else if (wbdata[22:12] == 991) begin 
      x02bai <= 32'b00111111101011000111110111010101;
      x02jyou <= 32'b00111110111010000111001010101000;
    end else if (wbdata[22:12] == 992) begin 
      x02bai <= 32'b00111111101011000110111101001111;
      x02jyou <= 32'b00111110111010000100101110000101;
    end else if (wbdata[22:12] == 993) begin 
      x02bai <= 32'b00111111101011000110000011001100;
      x02jyou <= 32'b00111110111010000010010001101101;
    end else if (wbdata[22:12] == 994) begin 
      x02bai <= 32'b00111111101011000101001001001011;
      x02jyou <= 32'b00111110111001111111110101011110;
    end else if (wbdata[22:12] == 995) begin 
      x02bai <= 32'b00111111101011000100001111001100;
      x02jyou <= 32'b00111110111001111101011001011000;
    end else if (wbdata[22:12] == 996) begin 
      x02bai <= 32'b00111111101011000011010101010000;
      x02jyou <= 32'b00111110111001111010111101011101;
    end else if (wbdata[22:12] == 997) begin 
      x02bai <= 32'b00111111101011000010011011010110;
      x02jyou <= 32'b00111110111001111000100001101011;
    end else if (wbdata[22:12] == 998) begin 
      x02bai <= 32'b00111111101011000001100001011111;
      x02jyou <= 32'b00111110111001110110000110000100;
    end else if (wbdata[22:12] == 999) begin 
      x02bai <= 32'b00111111101011000000100111101010;
      x02jyou <= 32'b00111110111001110011101010100110;
    end else if (wbdata[22:12] == 1000) begin 
      x02bai <= 32'b00111111101010111111101101110111;
      x02jyou <= 32'b00111110111001110001001111010000;
    end else if (wbdata[22:12] == 1001) begin 
      x02bai <= 32'b00111111101010111110110100000111;
      x02jyou <= 32'b00111110111001101110110100000110;
    end else if (wbdata[22:12] == 1002) begin 
      x02bai <= 32'b00111111101010111101111010011010;
      x02jyou <= 32'b00111110111001101100011001000111;
    end else if (wbdata[22:12] == 1003) begin 
      x02bai <= 32'b00111111101010111101000000101111;
      x02jyou <= 32'b00111110111001101001111110010000;
    end else if (wbdata[22:12] == 1004) begin 
      x02bai <= 32'b00111111101010111100000111000110;
      x02jyou <= 32'b00111110111001100111100011100010;
    end else if (wbdata[22:12] == 1005) begin 
      x02bai <= 32'b00111111101010111011001101100000;
      x02jyou <= 32'b00111110111001100101001001000000;
    end else if (wbdata[22:12] == 1006) begin 
      x02bai <= 32'b00111111101010111010010011111100;
      x02jyou <= 32'b00111110111001100010101110100110;
    end else if (wbdata[22:12] == 1007) begin 
      x02bai <= 32'b00111111101010111001011010011010;
      x02jyou <= 32'b00111110111001100000010100010101;
    end else if (wbdata[22:12] == 1008) begin 
      x02bai <= 32'b00111111101010111000100000111011;
      x02jyou <= 32'b00111110111001011101111010001111;
    end else if (wbdata[22:12] == 1009) begin 
      x02bai <= 32'b00111111101010110111100111011110;
      x02jyou <= 32'b00111110111001011011100000010001;
    end else if (wbdata[22:12] == 1010) begin 
      x02bai <= 32'b00111111101010110110101110000100;
      x02jyou <= 32'b00111110111001011001000110011111;
    end else if (wbdata[22:12] == 1011) begin 
      x02bai <= 32'b00111111101010110101110100101100;
      x02jyou <= 32'b00111110111001010110101100110101;
    end else if (wbdata[22:12] == 1012) begin 
      x02bai <= 32'b00111111101010110100111011010111;
      x02jyou <= 32'b00111110111001010100010011010111;
    end else if (wbdata[22:12] == 1013) begin 
      x02bai <= 32'b00111111101010110100000010000011;
      x02jyou <= 32'b00111110111001010001111001111111;
    end else if (wbdata[22:12] == 1014) begin 
      x02bai <= 32'b00111111101010110011001000110011;
      x02jyou <= 32'b00111110111001001111100000110100;
    end else if (wbdata[22:12] == 1015) begin 
      x02bai <= 32'b00111111101010110010001111100100;
      x02jyou <= 32'b00111110111001001101000111101111;
    end else if (wbdata[22:12] == 1016) begin 
      x02bai <= 32'b00111111101010110001010110011000;
      x02jyou <= 32'b00111110111001001010101110110110;
    end else if (wbdata[22:12] == 1017) begin 
      x02bai <= 32'b00111111101010110000011101001111;
      x02jyou <= 32'b00111110111001001000010110000111;
    end else if (wbdata[22:12] == 1018) begin 
      x02bai <= 32'b00111111101010101111100100001000;
      x02jyou <= 32'b00111110111001000101111101100010;
    end else if (wbdata[22:12] == 1019) begin 
      x02bai <= 32'b00111111101010101110101011000011;
      x02jyou <= 32'b00111110111001000011100101000101;
    end else if (wbdata[22:12] == 1020) begin 
      x02bai <= 32'b00111111101010101101110010000001;
      x02jyou <= 32'b00111110111001000001001100110011;
    end else if (wbdata[22:12] == 1021) begin 
      x02bai <= 32'b00111111101010101100111001000001;
      x02jyou <= 32'b00111110111000111110110100101001;
    end else if (wbdata[22:12] == 1022) begin 
      x02bai <= 32'b00111111101010101100000000000011;
      x02jyou <= 32'b00111110111000111100011100101000;
    end else if (wbdata[22:12] == 1023) begin 
      x02bai <= 32'b00111111101010101011000111001000;
      x02jyou <= 32'b00111110111000111010000100110010;
    end else if (wbdata[22:12] == 1024) begin 
      x02bai <= 32'b00111111101010101010001110001111;
      x02jyou <= 32'b00111110111000110111101101000101;
    end else if (wbdata[22:12] == 1025) begin 
      x02bai <= 32'b00111111101010101001010101011000;
      x02jyou <= 32'b00111110111000110101010101100000;
    end else if (wbdata[22:12] == 1026) begin 
      x02bai <= 32'b00111111101010101000011100100100;
      x02jyou <= 32'b00111110111000110010111110000110;
    end else if (wbdata[22:12] == 1027) begin 
      x02bai <= 32'b00111111101010100111100011110010;
      x02jyou <= 32'b00111110111000110000100110110101;
    end else if (wbdata[22:12] == 1028) begin 
      x02bai <= 32'b00111111101010100110101011000011;
      x02jyou <= 32'b00111110111000101110001111101111;
    end else if (wbdata[22:12] == 1029) begin 
      x02bai <= 32'b00111111101010100101110010010110;
      x02jyou <= 32'b00111110111000101011111000110001;
    end else if (wbdata[22:12] == 1030) begin 
      x02bai <= 32'b00111111101010100100111001101011;
      x02jyou <= 32'b00111110111000101001100001111100;
    end else if (wbdata[22:12] == 1031) begin 
      x02bai <= 32'b00111111101010100100000001000011;
      x02jyou <= 32'b00111110111000100111001011010010;
    end else if (wbdata[22:12] == 1032) begin 
      x02bai <= 32'b00111111101010100011001000011101;
      x02jyou <= 32'b00111110111000100100110100110001;
    end else if (wbdata[22:12] == 1033) begin 
      x02bai <= 32'b00111111101010100010001111111001;
      x02jyou <= 32'b00111110111000100010011110011000;
    end else if (wbdata[22:12] == 1034) begin 
      x02bai <= 32'b00111111101010100001010111011000;
      x02jyou <= 32'b00111110111000100000001000001001;
    end else if (wbdata[22:12] == 1035) begin 
      x02bai <= 32'b00111111101010100000011110111001;
      x02jyou <= 32'b00111110111000011101110010000100;
    end else if (wbdata[22:12] == 1036) begin 
      x02bai <= 32'b00111111101010011111100110011100;
      x02jyou <= 32'b00111110111000011011011100000111;
    end else if (wbdata[22:12] == 1037) begin 
      x02bai <= 32'b00111111101010011110101110000010;
      x02jyou <= 32'b00111110111000011001000110010101;
    end else if (wbdata[22:12] == 1038) begin 
      x02bai <= 32'b00111111101010011101110101101010;
      x02jyou <= 32'b00111110111000010110110000101011;
    end else if (wbdata[22:12] == 1039) begin 
      x02bai <= 32'b00111111101010011100111101010100;
      x02jyou <= 32'b00111110111000010100011011001010;
    end else if (wbdata[22:12] == 1040) begin 
      x02bai <= 32'b00111111101010011100000101000001;
      x02jyou <= 32'b00111110111000010010000101110011;
    end else if (wbdata[22:12] == 1041) begin 
      x02bai <= 32'b00111111101010011011001100110000;
      x02jyou <= 32'b00111110111000001111110000100110;
    end else if (wbdata[22:12] == 1042) begin 
      x02bai <= 32'b00111111101010011010010100100010;
      x02jyou <= 32'b00111110111000001101011011100011;
    end else if (wbdata[22:12] == 1043) begin 
      x02bai <= 32'b00111111101010011001011100010101;
      x02jyou <= 32'b00111110111000001011000110100110;
    end else if (wbdata[22:12] == 1044) begin 
      x02bai <= 32'b00111111101010011000100100001100;
      x02jyou <= 32'b00111110111000001000110001110110;
    end else if (wbdata[22:12] == 1045) begin 
      x02bai <= 32'b00111111101010010111101100000100;
      x02jyou <= 32'b00111110111000000110011101001101;
    end else if (wbdata[22:12] == 1046) begin 
      x02bai <= 32'b00111111101010010110110011111111;
      x02jyou <= 32'b00111110111000000100001000101110;
    end else if (wbdata[22:12] == 1047) begin 
      x02bai <= 32'b00111111101010010101111011111100;
      x02jyou <= 32'b00111110111000000001110100011000;
    end else if (wbdata[22:12] == 1048) begin 
      x02bai <= 32'b00111111101010010101000011111011;
      x02jyou <= 32'b00111110110111111111100000001010;
    end else if (wbdata[22:12] == 1049) begin 
      x02bai <= 32'b00111111101010010100001011111101;
      x02jyou <= 32'b00111110110111111101001100000111;
    end else if (wbdata[22:12] == 1050) begin 
      x02bai <= 32'b00111111101010010011010100000001;
      x02jyou <= 32'b00111110110111111010111000001101;
    end else if (wbdata[22:12] == 1051) begin 
      x02bai <= 32'b00111111101010010010011100000111;
      x02jyou <= 32'b00111110110111111000100100011010;
    end else if (wbdata[22:12] == 1052) begin 
      x02bai <= 32'b00111111101010010001100100001111;
      x02jyou <= 32'b00111110110111110110010000110001;
    end else if (wbdata[22:12] == 1053) begin 
      x02bai <= 32'b00111111101010010000101100011010;
      x02jyou <= 32'b00111110110111110011111101010010;
    end else if (wbdata[22:12] == 1054) begin 
      x02bai <= 32'b00111111101010001111110100101000;
      x02jyou <= 32'b00111110110111110001101001111110;
    end else if (wbdata[22:12] == 1055) begin 
      x02bai <= 32'b00111111101010001110111100110111;
      x02jyou <= 32'b00111110110111101111010110101111;
    end else if (wbdata[22:12] == 1056) begin 
      x02bai <= 32'b00111111101010001110000101001001;
      x02jyou <= 32'b00111110110111101101000011101100;
    end else if (wbdata[22:12] == 1057) begin 
      x02bai <= 32'b00111111101010001101001101011101;
      x02jyou <= 32'b00111110110111101010110000110001;
    end else if (wbdata[22:12] == 1058) begin 
      x02bai <= 32'b00111111101010001100010101110011;
      x02jyou <= 32'b00111110110111101000011101111110;
    end else if (wbdata[22:12] == 1059) begin 
      x02bai <= 32'b00111111101010001011011110001100;
      x02jyou <= 32'b00111110110111100110001011010111;
    end else if (wbdata[22:12] == 1060) begin 
      x02bai <= 32'b00111111101010001010100110100111;
      x02jyou <= 32'b00111110110111100011111000110111;
    end else if (wbdata[22:12] == 1061) begin 
      x02bai <= 32'b00111111101010001001101111000100;
      x02jyou <= 32'b00111110110111100001100110100000;
    end else if (wbdata[22:12] == 1062) begin 
      x02bai <= 32'b00111111101010001000110111100100;
      x02jyou <= 32'b00111110110111011111010100010100;
    end else if (wbdata[22:12] == 1063) begin 
      x02bai <= 32'b00111111101010001000000000000110;
      x02jyou <= 32'b00111110110111011101000010010000;
    end else if (wbdata[22:12] == 1064) begin 
      x02bai <= 32'b00111111101010000111001000101010;
      x02jyou <= 32'b00111110110111011010110000010100;
    end else if (wbdata[22:12] == 1065) begin 
      x02bai <= 32'b00111111101010000110010001010000;
      x02jyou <= 32'b00111110110111011000011110100001;
    end else if (wbdata[22:12] == 1066) begin 
      x02bai <= 32'b00111111101010000101011001111001;
      x02jyou <= 32'b00111110110111010110001100111000;
    end else if (wbdata[22:12] == 1067) begin 
      x02bai <= 32'b00111111101010000100100010100100;
      x02jyou <= 32'b00111110110111010011111011011000;
    end else if (wbdata[22:12] == 1068) begin 
      x02bai <= 32'b00111111101010000011101011010001;
      x02jyou <= 32'b00111110110111010001101010000000;
    end else if (wbdata[22:12] == 1069) begin 
      x02bai <= 32'b00111111101010000010110100000000;
      x02jyou <= 32'b00111110110111001111011000110000;
    end else if (wbdata[22:12] == 1070) begin 
      x02bai <= 32'b00111111101010000001111100110010;
      x02jyou <= 32'b00111110110111001101000111101011;
    end else if (wbdata[22:12] == 1071) begin 
      x02bai <= 32'b00111111101010000001000101100110;
      x02jyou <= 32'b00111110110111001010110110101110;
    end else if (wbdata[22:12] == 1072) begin 
      x02bai <= 32'b00111111101010000000001110011100;
      x02jyou <= 32'b00111110110111001000100101111010;
    end else if (wbdata[22:12] == 1073) begin 
      x02bai <= 32'b00111111101001111111010111010101;
      x02jyou <= 32'b00111110110111000110010101010000;
    end else if (wbdata[22:12] == 1074) begin 
      x02bai <= 32'b00111111101001111110100000010000;
      x02jyou <= 32'b00111110110111000100000100101110;
    end else if (wbdata[22:12] == 1075) begin 
      x02bai <= 32'b00111111101001111101101001001101;
      x02jyou <= 32'b00111110110111000001110100010101;
    end else if (wbdata[22:12] == 1076) begin 
      x02bai <= 32'b00111111101001111100110010001100;
      x02jyou <= 32'b00111110110110111111100100000100;
    end else if (wbdata[22:12] == 1077) begin 
      x02bai <= 32'b00111111101001111011111011001110;
      x02jyou <= 32'b00111110110110111101010011111110;
    end else if (wbdata[22:12] == 1078) begin 
      x02bai <= 32'b00111111101001111011000100010001;
      x02jyou <= 32'b00111110110110111011000011111101;
    end else if (wbdata[22:12] == 1079) begin 
      x02bai <= 32'b00111111101001111010001101010111;
      x02jyou <= 32'b00111110110110111000110100000111;
    end else if (wbdata[22:12] == 1080) begin 
      x02bai <= 32'b00111111101001111001010110100000;
      x02jyou <= 32'b00111110110110110110100100011100;
    end else if (wbdata[22:12] == 1081) begin 
      x02bai <= 32'b00111111101001111000011111101010;
      x02jyou <= 32'b00111110110110110100010100110111;
    end else if (wbdata[22:12] == 1082) begin 
      x02bai <= 32'b00111111101001110111101000110111;
      x02jyou <= 32'b00111110110110110010000101011100;
    end else if (wbdata[22:12] == 1083) begin 
      x02bai <= 32'b00111111101001110110110010000110;
      x02jyou <= 32'b00111110110110101111110110001010;
    end else if (wbdata[22:12] == 1084) begin 
      x02bai <= 32'b00111111101001110101111011010111;
      x02jyou <= 32'b00111110110110101101100110111111;
    end else if (wbdata[22:12] == 1085) begin 
      x02bai <= 32'b00111111101001110101000100101011;
      x02jyou <= 32'b00111110110110101011011000000000;
    end else if (wbdata[22:12] == 1086) begin 
      x02bai <= 32'b00111111101001110100001110000001;
      x02jyou <= 32'b00111110110110101001001001001000;
    end else if (wbdata[22:12] == 1087) begin 
      x02bai <= 32'b00111111101001110011010111011001;
      x02jyou <= 32'b00111110110110100110111010011001;
    end else if (wbdata[22:12] == 1088) begin 
      x02bai <= 32'b00111111101001110010100000110011;
      x02jyou <= 32'b00111110110110100100101011110010;
    end else if (wbdata[22:12] == 1089) begin 
      x02bai <= 32'b00111111101001110001101010001111;
      x02jyou <= 32'b00111110110110100010011101010011;
    end else if (wbdata[22:12] == 1090) begin 
      x02bai <= 32'b00111111101001110000110011101110;
      x02jyou <= 32'b00111110110110100000001110111110;
    end else if (wbdata[22:12] == 1091) begin 
      x02bai <= 32'b00111111101001101111111101001111;
      x02jyou <= 32'b00111110110110011110000000110010;
    end else if (wbdata[22:12] == 1092) begin 
      x02bai <= 32'b00111111101001101111000110110010;
      x02jyou <= 32'b00111110110110011011110010101110;
    end else if (wbdata[22:12] == 1093) begin 
      x02bai <= 32'b00111111101001101110010000010111;
      x02jyou <= 32'b00111110110110011001100100110010;
    end else if (wbdata[22:12] == 1094) begin 
      x02bai <= 32'b00111111101001101101011001111111;
      x02jyou <= 32'b00111110110110010111010111000001;
    end else if (wbdata[22:12] == 1095) begin 
      x02bai <= 32'b00111111101001101100100011101001;
      x02jyou <= 32'b00111110110110010101001001011000;
    end else if (wbdata[22:12] == 1096) begin 
      x02bai <= 32'b00111111101001101011101101010100;
      x02jyou <= 32'b00111110110110010010111011110100;
    end else if (wbdata[22:12] == 1097) begin 
      x02bai <= 32'b00111111101001101010110111000011;
      x02jyou <= 32'b00111110110110010000101110011110;
    end else if (wbdata[22:12] == 1098) begin 
      x02bai <= 32'b00111111101001101010000000110011;
      x02jyou <= 32'b00111110110110001110100001001101;
    end else if (wbdata[22:12] == 1099) begin 
      x02bai <= 32'b00111111101001101001001010100110;
      x02jyou <= 32'b00111110110110001100010100000111;
    end else if (wbdata[22:12] == 1100) begin 
      x02bai <= 32'b00111111101001101000010100011010;
      x02jyou <= 32'b00111110110110001010000111000110;
    end else if (wbdata[22:12] == 1101) begin 
      x02bai <= 32'b00111111101001100111011110010001;
      x02jyou <= 32'b00111110110110000111111010010000;
    end else if (wbdata[22:12] == 1102) begin 
      x02bai <= 32'b00111111101001100110101000001011;
      x02jyou <= 32'b00111110110110000101101101100100;
    end else if (wbdata[22:12] == 1103) begin 
      x02bai <= 32'b00111111101001100101110010000110;
      x02jyou <= 32'b00111110110110000011100000111110;
    end else if (wbdata[22:12] == 1104) begin 
      x02bai <= 32'b00111111101001100100111100000100;
      x02jyou <= 32'b00111110110110000001010100100011;
    end else if (wbdata[22:12] == 1105) begin 
      x02bai <= 32'b00111111101001100100000110000011;
      x02jyou <= 32'b00111110110101111111001000001101;
    end else if (wbdata[22:12] == 1106) begin 
      x02bai <= 32'b00111111101001100011010000000101;
      x02jyou <= 32'b00111110110101111100111100000010;
    end else if (wbdata[22:12] == 1107) begin 
      x02bai <= 32'b00111111101001100010011010001001;
      x02jyou <= 32'b00111110110101111010101111111111;
    end else if (wbdata[22:12] == 1108) begin 
      x02bai <= 32'b00111111101001100001100100010000;
      x02jyou <= 32'b00111110110101111000100100000110;
    end else if (wbdata[22:12] == 1109) begin 
      x02bai <= 32'b00111111101001100000101110011000;
      x02jyou <= 32'b00111110110101110110011000010011;
    end else if (wbdata[22:12] == 1110) begin 
      x02bai <= 32'b00111111101001011111111000100011;
      x02jyou <= 32'b00111110110101110100001100101011;
    end else if (wbdata[22:12] == 1111) begin 
      x02bai <= 32'b00111111101001011111000010110000;
      x02jyou <= 32'b00111110110101110010000001001010;
    end else if (wbdata[22:12] == 1112) begin 
      x02bai <= 32'b00111111101001011110001100111111;
      x02jyou <= 32'b00111110110101101111110101110010;
    end else if (wbdata[22:12] == 1113) begin 
      x02bai <= 32'b00111111101001011101010111010000;
      x02jyou <= 32'b00111110110101101101101010100001;
    end else if (wbdata[22:12] == 1114) begin 
      x02bai <= 32'b00111111101001011100100001100100;
      x02jyou <= 32'b00111110110101101011011111011100;
    end else if (wbdata[22:12] == 1115) begin 
      x02bai <= 32'b00111111101001011011101011111001;
      x02jyou <= 32'b00111110110101101001010100011011;
    end else if (wbdata[22:12] == 1116) begin 
      x02bai <= 32'b00111111101001011010110110010001;
      x02jyou <= 32'b00111110110101100111001001100101;
    end else if (wbdata[22:12] == 1117) begin 
      x02bai <= 32'b00111111101001011010000000101011;
      x02jyou <= 32'b00111110110101100100111110110111;
    end else if (wbdata[22:12] == 1118) begin 
      x02bai <= 32'b00111111101001011001001011000111;
      x02jyou <= 32'b00111110110101100010110100010001;
    end else if (wbdata[22:12] == 1119) begin 
      x02bai <= 32'b00111111101001011000010101100101;
      x02jyou <= 32'b00111110110101100000101001110011;
    end else if (wbdata[22:12] == 1120) begin 
      x02bai <= 32'b00111111101001010111100000000110;
      x02jyou <= 32'b00111110110101011110011111100000;
    end else if (wbdata[22:12] == 1121) begin 
      x02bai <= 32'b00111111101001010110101010101000;
      x02jyou <= 32'b00111110110101011100010101010010;
    end else if (wbdata[22:12] == 1122) begin 
      x02bai <= 32'b00111111101001010101110101001101;
      x02jyou <= 32'b00111110110101011010001011001111;
    end else if (wbdata[22:12] == 1123) begin 
      x02bai <= 32'b00111111101001010100111111110100;
      x02jyou <= 32'b00111110110101011000000001010011;
    end else if (wbdata[22:12] == 1124) begin 
      x02bai <= 32'b00111111101001010100001010011101;
      x02jyou <= 32'b00111110110101010101110111011111;
    end else if (wbdata[22:12] == 1125) begin 
      x02bai <= 32'b00111111101001010011010101001000;
      x02jyou <= 32'b00111110110101010011101101110100;
    end else if (wbdata[22:12] == 1126) begin 
      x02bai <= 32'b00111111101001010010011111110110;
      x02jyou <= 32'b00111110110101010001100100010011;
    end else if (wbdata[22:12] == 1127) begin 
      x02bai <= 32'b00111111101001010001101010100101;
      x02jyou <= 32'b00111110110101001111011010110111;
    end else if (wbdata[22:12] == 1128) begin 
      x02bai <= 32'b00111111101001010000110101010111;
      x02jyou <= 32'b00111110110101001101010001100110;
    end else if (wbdata[22:12] == 1129) begin 
      x02bai <= 32'b00111111101001010000000000001011;
      x02jyou <= 32'b00111110110101001011001000011100;
    end else if (wbdata[22:12] == 1130) begin 
      x02bai <= 32'b00111111101001001111001011000001;
      x02jyou <= 32'b00111110110101001000111111011011;
    end else if (wbdata[22:12] == 1131) begin 
      x02bai <= 32'b00111111101001001110010101111001;
      x02jyou <= 32'b00111110110101000110110110100001;
    end else if (wbdata[22:12] == 1132) begin 
      x02bai <= 32'b00111111101001001101100000110011;
      x02jyou <= 32'b00111110110101000100101101110000;
    end else if (wbdata[22:12] == 1133) begin 
      x02bai <= 32'b00111111101001001100101011101111;
      x02jyou <= 32'b00111110110101000010100101000110;
    end else if (wbdata[22:12] == 1134) begin 
      x02bai <= 32'b00111111101001001011110110101110;
      x02jyou <= 32'b00111110110101000000011100100111;
    end else if (wbdata[22:12] == 1135) begin 
      x02bai <= 32'b00111111101001001011000001101110;
      x02jyou <= 32'b00111110110100111110010100001101;
    end else if (wbdata[22:12] == 1136) begin 
      x02bai <= 32'b00111111101001001010001100110001;
      x02jyou <= 32'b00111110110100111100001011111110;
    end else if (wbdata[22:12] == 1137) begin 
      x02bai <= 32'b00111111101001001001010111110110;
      x02jyou <= 32'b00111110110100111010000011110110;
    end else if (wbdata[22:12] == 1138) begin 
      x02bai <= 32'b00111111101001001000100010111101;
      x02jyou <= 32'b00111110110100110111111011110110;
    end else if (wbdata[22:12] == 1139) begin 
      x02bai <= 32'b00111111101001000111101110000110;
      x02jyou <= 32'b00111110110100110101110011111111;
    end else if (wbdata[22:12] == 1140) begin 
      x02bai <= 32'b00111111101001000110111001010001;
      x02jyou <= 32'b00111110110100110011101100001111;
    end else if (wbdata[22:12] == 1141) begin 
      x02bai <= 32'b00111111101001000110000100011111;
      x02jyou <= 32'b00111110110100110001100100101001;
    end else if (wbdata[22:12] == 1142) begin 
      x02bai <= 32'b00111111101001000101001111101110;
      x02jyou <= 32'b00111110110100101111011101001001;
    end else if (wbdata[22:12] == 1143) begin 
      x02bai <= 32'b00111111101001000100011011000000;
      x02jyou <= 32'b00111110110100101101010101110011;
    end else if (wbdata[22:12] == 1144) begin 
      x02bai <= 32'b00111111101001000011100110010011;
      x02jyou <= 32'b00111110110100101011001110100011;
    end else if (wbdata[22:12] == 1145) begin 
      x02bai <= 32'b00111111101001000010110001101001;
      x02jyou <= 32'b00111110110100101001000111011100;
    end else if (wbdata[22:12] == 1146) begin 
      x02bai <= 32'b00111111101001000001111101000001;
      x02jyou <= 32'b00111110110100100111000000011110;
    end else if (wbdata[22:12] == 1147) begin 
      x02bai <= 32'b00111111101001000001001000011011;
      x02jyou <= 32'b00111110110100100100111001101000;
    end else if (wbdata[22:12] == 1148) begin 
      x02bai <= 32'b00111111101001000000010011110111;
      x02jyou <= 32'b00111110110100100010110010111001;
    end else if (wbdata[22:12] == 1149) begin 
      x02bai <= 32'b00111111101000111111011111010110;
      x02jyou <= 32'b00111110110100100000101100010101;
    end else if (wbdata[22:12] == 1150) begin 
      x02bai <= 32'b00111111101000111110101010110110;
      x02jyou <= 32'b00111110110100011110100101110110;
    end else if (wbdata[22:12] == 1151) begin 
      x02bai <= 32'b00111111101000111101110110011000;
      x02jyou <= 32'b00111110110100011100011111011111;
    end else if (wbdata[22:12] == 1152) begin 
      x02bai <= 32'b00111111101000111101000001111101;
      x02jyou <= 32'b00111110110100011010011001010010;
    end else if (wbdata[22:12] == 1153) begin 
      x02bai <= 32'b00111111101000111100001101100100;
      x02jyou <= 32'b00111110110100011000010011001101;
    end else if (wbdata[22:12] == 1154) begin 
      x02bai <= 32'b00111111101000111011011001001100;
      x02jyou <= 32'b00111110110100010110001101001101;
    end else if (wbdata[22:12] == 1155) begin 
      x02bai <= 32'b00111111101000111010100100110111;
      x02jyou <= 32'b00111110110100010100000111011000;
    end else if (wbdata[22:12] == 1156) begin 
      x02bai <= 32'b00111111101000111001110000100100;
      x02jyou <= 32'b00111110110100010010000001101010;
    end else if (wbdata[22:12] == 1157) begin 
      x02bai <= 32'b00111111101000111000111100010011;
      x02jyou <= 32'b00111110110100001111111100000100;
    end else if (wbdata[22:12] == 1158) begin 
      x02bai <= 32'b00111111101000111000001000000100;
      x02jyou <= 32'b00111110110100001101110110100110;
    end else if (wbdata[22:12] == 1159) begin 
      x02bai <= 32'b00111111101000110111010011111000;
      x02jyou <= 32'b00111110110100001011110001010011;
    end else if (wbdata[22:12] == 1160) begin 
      x02bai <= 32'b00111111101000110110011111101101;
      x02jyou <= 32'b00111110110100001001101100000100;
    end else if (wbdata[22:12] == 1161) begin 
      x02bai <= 32'b00111111101000110101101011100100;
      x02jyou <= 32'b00111110110100000111100110111101;
    end else if (wbdata[22:12] == 1162) begin 
      x02bai <= 32'b00111111101000110100110111011110;
      x02jyou <= 32'b00111110110100000101100010000001;
    end else if (wbdata[22:12] == 1163) begin 
      x02bai <= 32'b00111111101000110100000011011001;
      x02jyou <= 32'b00111110110100000011011101001010;
    end else if (wbdata[22:12] == 1164) begin 
      x02bai <= 32'b00111111101000110011001111010111;
      x02jyou <= 32'b00111110110100000001011000011101;
    end else if (wbdata[22:12] == 1165) begin 
      x02bai <= 32'b00111111101000110010011011010110;
      x02jyou <= 32'b00111110110011111111010011110101;
    end else if (wbdata[22:12] == 1166) begin 
      x02bai <= 32'b00111111101000110001100111011000;
      x02jyou <= 32'b00111110110011111101001111010111;
    end else if (wbdata[22:12] == 1167) begin 
      x02bai <= 32'b00111111101000110000110011011100;
      x02jyou <= 32'b00111110110011111011001011000010;
    end else if (wbdata[22:12] == 1168) begin 
      x02bai <= 32'b00111111101000101111111111100010;
      x02jyou <= 32'b00111110110011111001000110110100;
    end else if (wbdata[22:12] == 1169) begin 
      x02bai <= 32'b00111111101000101111001011101010;
      x02jyou <= 32'b00111110110011110111000010101101;
    end else if (wbdata[22:12] == 1170) begin 
      x02bai <= 32'b00111111101000101110010111110100;
      x02jyou <= 32'b00111110110011110100111110101111;
    end else if (wbdata[22:12] == 1171) begin 
      x02bai <= 32'b00111111101000101101100100000000;
      x02jyou <= 32'b00111110110011110010111010111000;
    end else if (wbdata[22:12] == 1172) begin 
      x02bai <= 32'b00111111101000101100110000001110;
      x02jyou <= 32'b00111110110011110000110111001001;
    end else if (wbdata[22:12] == 1173) begin 
      x02bai <= 32'b00111111101000101011111100011110;
      x02jyou <= 32'b00111110110011101110110011100001;
    end else if (wbdata[22:12] == 1174) begin 
      x02bai <= 32'b00111111101000101011001000110000;
      x02jyou <= 32'b00111110110011101100110000000010;
    end else if (wbdata[22:12] == 1175) begin 
      x02bai <= 32'b00111111101000101010010101000100;
      x02jyou <= 32'b00111110110011101010101100101010;
    end else if (wbdata[22:12] == 1176) begin 
      x02bai <= 32'b00111111101000101001100001011011;
      x02jyou <= 32'b00111110110011101000101001011100;
    end else if (wbdata[22:12] == 1177) begin 
      x02bai <= 32'b00111111101000101000101101110011;
      x02jyou <= 32'b00111110110011100110100110010011;
    end else if (wbdata[22:12] == 1178) begin 
      x02bai <= 32'b00111111101000100111111010001110;
      x02jyou <= 32'b00111110110011100100100011010101;
    end else if (wbdata[22:12] == 1179) begin 
      x02bai <= 32'b00111111101000100111000110101010;
      x02jyou <= 32'b00111110110011100010100000011011;
    end else if (wbdata[22:12] == 1180) begin 
      x02bai <= 32'b00111111101000100110010011001001;
      x02jyou <= 32'b00111110110011100000011101101100;
    end else if (wbdata[22:12] == 1181) begin 
      x02bai <= 32'b00111111101000100101011111101001;
      x02jyou <= 32'b00111110110011011110011011000010;
    end else if (wbdata[22:12] == 1182) begin 
      x02bai <= 32'b00111111101000100100101100001100;
      x02jyou <= 32'b00111110110011011100011000100010;
    end else if (wbdata[22:12] == 1183) begin 
      x02bai <= 32'b00111111101000100011111000110000;
      x02jyou <= 32'b00111110110011011010010110001000;
    end else if (wbdata[22:12] == 1184) begin 
      x02bai <= 32'b00111111101000100011000101010111;
      x02jyou <= 32'b00111110110011011000010011110111;
    end else if (wbdata[22:12] == 1185) begin 
      x02bai <= 32'b00111111101000100010010010000000;
      x02jyou <= 32'b00111110110011010110010001101110;
    end else if (wbdata[22:12] == 1186) begin 
      x02bai <= 32'b00111111101000100001011110101010;
      x02jyou <= 32'b00111110110011010100001111101011;
    end else if (wbdata[22:12] == 1187) begin 
      x02bai <= 32'b00111111101000100000101011010111;
      x02jyou <= 32'b00111110110011010010001101110001;
    end else if (wbdata[22:12] == 1188) begin 
      x02bai <= 32'b00111111101000011111111000000110;
      x02jyou <= 32'b00111110110011010000001011111111;
    end else if (wbdata[22:12] == 1189) begin 
      x02bai <= 32'b00111111101000011111000100110111;
      x02jyou <= 32'b00111110110011001110001010010101;
    end else if (wbdata[22:12] == 1190) begin 
      x02bai <= 32'b00111111101000011110010001101010;
      x02jyou <= 32'b00111110110011001100001000110010;
    end else if (wbdata[22:12] == 1191) begin 
      x02bai <= 32'b00111111101000011101011110011111;
      x02jyou <= 32'b00111110110011001010000111010111;
    end else if (wbdata[22:12] == 1192) begin 
      x02bai <= 32'b00111111101000011100101011010101;
      x02jyou <= 32'b00111110110011001000000110000001;
    end else if (wbdata[22:12] == 1193) begin 
      x02bai <= 32'b00111111101000011011111000001110;
      x02jyou <= 32'b00111110110011000110000100110101;
    end else if (wbdata[22:12] == 1194) begin 
      x02bai <= 32'b00111111101000011011000101001001;
      x02jyou <= 32'b00111110110011000100000011110001;
    end else if (wbdata[22:12] == 1195) begin 
      x02bai <= 32'b00111111101000011010010010000110;
      x02jyou <= 32'b00111110110011000010000010110101;
    end else if (wbdata[22:12] == 1196) begin 
      x02bai <= 32'b00111111101000011001011111000101;
      x02jyou <= 32'b00111110110011000000000010000000;
    end else if (wbdata[22:12] == 1197) begin 
      x02bai <= 32'b00111111101000011000101100000110;
      x02jyou <= 32'b00111110110010111110000001010010;
    end else if (wbdata[22:12] == 1198) begin 
      x02bai <= 32'b00111111101000010111111001001001;
      x02jyou <= 32'b00111110110010111100000000101100;
    end else if (wbdata[22:12] == 1199) begin 
      x02bai <= 32'b00111111101000010111000110001110;
      x02jyou <= 32'b00111110110010111010000000001110;
    end else if (wbdata[22:12] == 1200) begin 
      x02bai <= 32'b00111111101000010110010011010101;
      x02jyou <= 32'b00111110110010110111111111110111;
    end else if (wbdata[22:12] == 1201) begin 
      x02bai <= 32'b00111111101000010101100000011110;
      x02jyou <= 32'b00111110110010110101111111101000;
    end else if (wbdata[22:12] == 1202) begin 
      x02bai <= 32'b00111111101000010100101101101001;
      x02jyou <= 32'b00111110110010110011111111100001;
    end else if (wbdata[22:12] == 1203) begin 
      x02bai <= 32'b00111111101000010011111010110110;
      x02jyou <= 32'b00111110110010110001111111100001;
    end else if (wbdata[22:12] == 1204) begin 
      x02bai <= 32'b00111111101000010011001000000101;
      x02jyou <= 32'b00111110110010101111111111101000;
    end else if (wbdata[22:12] == 1205) begin 
      x02bai <= 32'b00111111101000010010010101010110;
      x02jyou <= 32'b00111110110010101101111111110111;
    end else if (wbdata[22:12] == 1206) begin 
      x02bai <= 32'b00111111101000010001100010101001;
      x02jyou <= 32'b00111110110010101100000000001110;
    end else if (wbdata[22:12] == 1207) begin 
      x02bai <= 32'b00111111101000010000101111111110;
      x02jyou <= 32'b00111110110010101010000000101100;
    end else if (wbdata[22:12] == 1208) begin 
      x02bai <= 32'b00111111101000001111111101010101;
      x02jyou <= 32'b00111110110010101000000001010010;
    end else if (wbdata[22:12] == 1209) begin 
      x02bai <= 32'b00111111101000001111001010101110;
      x02jyou <= 32'b00111110110010100110000001111111;
    end else if (wbdata[22:12] == 1210) begin 
      x02bai <= 32'b00111111101000001110011000001001;
      x02jyou <= 32'b00111110110010100100000010110100;
    end else if (wbdata[22:12] == 1211) begin 
      x02bai <= 32'b00111111101000001101100101100110;
      x02jyou <= 32'b00111110110010100010000011110000;
    end else if (wbdata[22:12] == 1212) begin 
      x02bai <= 32'b00111111101000001100110011000101;
      x02jyou <= 32'b00111110110010100000000100110100;
    end else if (wbdata[22:12] == 1213) begin 
      x02bai <= 32'b00111111101000001100000000100110;
      x02jyou <= 32'b00111110110010011110000101111111;
    end else if (wbdata[22:12] == 1214) begin 
      x02bai <= 32'b00111111101000001011001110001001;
      x02jyou <= 32'b00111110110010011100000111010010;
    end else if (wbdata[22:12] == 1215) begin 
      x02bai <= 32'b00111111101000001010011011101110;
      x02jyou <= 32'b00111110110010011010001000101101;
    end else if (wbdata[22:12] == 1216) begin 
      x02bai <= 32'b00111111101000001001101001010101;
      x02jyou <= 32'b00111110110010011000001010001111;
    end else if (wbdata[22:12] == 1217) begin 
      x02bai <= 32'b00111111101000001000110110111101;
      x02jyou <= 32'b00111110110010010110001011110101;
    end else if (wbdata[22:12] == 1218) begin 
      x02bai <= 32'b00111111101000001000000100101000;
      x02jyou <= 32'b00111110110010010100001101100110;
    end else if (wbdata[22:12] == 1219) begin 
      x02bai <= 32'b00111111101000000111010010010101;
      x02jyou <= 32'b00111110110010010010001111011111;
    end else if (wbdata[22:12] == 1220) begin 
      x02bai <= 32'b00111111101000000110100000000100;
      x02jyou <= 32'b00111110110010010000010001011111;
    end else if (wbdata[22:12] == 1221) begin 
      x02bai <= 32'b00111111101000000101101101110100;
      x02jyou <= 32'b00111110110010001110010011100011;
    end else if (wbdata[22:12] == 1222) begin 
      x02bai <= 32'b00111111101000000100111011100111;
      x02jyou <= 32'b00111110110010001100010101110010;
    end else if (wbdata[22:12] == 1223) begin 
      x02bai <= 32'b00111111101000000100001001011100;
      x02jyou <= 32'b00111110110010001010011000001000;
    end else if (wbdata[22:12] == 1224) begin 
      x02bai <= 32'b00111111101000000011010111010010;
      x02jyou <= 32'b00111110110010001000011010100100;
    end else if (wbdata[22:12] == 1225) begin 
      x02bai <= 32'b00111111101000000010100101001011;
      x02jyou <= 32'b00111110110010000110011101001001;
    end else if (wbdata[22:12] == 1226) begin 
      x02bai <= 32'b00111111101000000001110011000101;
      x02jyou <= 32'b00111110110010000100011111110011;
    end else if (wbdata[22:12] == 1227) begin 
      x02bai <= 32'b00111111101000000001000001000010;
      x02jyou <= 32'b00111110110010000010100010100111;
    end else if (wbdata[22:12] == 1228) begin 
      x02bai <= 32'b00111111101000000000001111000000;
      x02jyou <= 32'b00111110110010000000100101100000;
    end else if (wbdata[22:12] == 1229) begin 
      x02bai <= 32'b00111111100111111111011101000001;
      x02jyou <= 32'b00111110110001111110101000100011;
    end else if (wbdata[22:12] == 1230) begin 
      x02bai <= 32'b00111111100111111110101011000011;
      x02jyou <= 32'b00111110110001111100101011101011;
    end else if (wbdata[22:12] == 1231) begin 
      x02bai <= 32'b00111111100111111101111001000111;
      x02jyou <= 32'b00111110110001111010101110111010;
    end else if (wbdata[22:12] == 1232) begin 
      x02bai <= 32'b00111111100111111101000111001110;
      x02jyou <= 32'b00111110110001111000110010010100;
    end else if (wbdata[22:12] == 1233) begin 
      x02bai <= 32'b00111111100111111100010101010110;
      x02jyou <= 32'b00111110110001110110110101110010;
    end else if (wbdata[22:12] == 1234) begin 
      x02bai <= 32'b00111111100111111011100011100000;
      x02jyou <= 32'b00111110110001110100111001011000;
    end else if (wbdata[22:12] == 1235) begin 
      x02bai <= 32'b00111111100111111010110001101100;
      x02jyou <= 32'b00111110110001110010111101000101;
    end else if (wbdata[22:12] == 1236) begin 
      x02bai <= 32'b00111111100111111001111111111010;
      x02jyou <= 32'b00111110110001110001000000111001;
    end else if (wbdata[22:12] == 1237) begin 
      x02bai <= 32'b00111111100111111001001110001010;
      x02jyou <= 32'b00111110110001101111000100110101;
    end else if (wbdata[22:12] == 1238) begin 
      x02bai <= 32'b00111111100111111000011100011100;
      x02jyou <= 32'b00111110110001101101001000111000;
    end else if (wbdata[22:12] == 1239) begin 
      x02bai <= 32'b00111111100111110111101010110000;
      x02jyou <= 32'b00111110110001101011001101000011;
    end else if (wbdata[22:12] == 1240) begin 
      x02bai <= 32'b00111111100111110110111001000101;
      x02jyou <= 32'b00111110110001101001010001010010;
    end else if (wbdata[22:12] == 1241) begin 
      x02bai <= 32'b00111111100111110110000111011101;
      x02jyou <= 32'b00111110110001100111010101101100;
    end else if (wbdata[22:12] == 1242) begin 
      x02bai <= 32'b00111111100111110101010101110111;
      x02jyou <= 32'b00111110110001100101011010001101;
    end else if (wbdata[22:12] == 1243) begin 
      x02bai <= 32'b00111111100111110100100100010010;
      x02jyou <= 32'b00111110110001100011011110110010;
    end else if (wbdata[22:12] == 1244) begin 
      x02bai <= 32'b00111111100111110011110010110000;
      x02jyou <= 32'b00111110110001100001100011100010;
    end else if (wbdata[22:12] == 1245) begin 
      x02bai <= 32'b00111111100111110011000001001111;
      x02jyou <= 32'b00111110110001011111101000010110;
    end else if (wbdata[22:12] == 1246) begin 
      x02bai <= 32'b00111111100111110010001111110001;
      x02jyou <= 32'b00111110110001011101101101010101;
    end else if (wbdata[22:12] == 1247) begin 
      x02bai <= 32'b00111111100111110001011110010100;
      x02jyou <= 32'b00111110110001011011110010011000;
    end else if (wbdata[22:12] == 1248) begin 
      x02bai <= 32'b00111111100111110000101100111001;
      x02jyou <= 32'b00111110110001011001110111100011;
    end else if (wbdata[22:12] == 1249) begin 
      x02bai <= 32'b00111111100111101111111011100000;
      x02jyou <= 32'b00111110110001010111111100110101;
    end else if (wbdata[22:12] == 1250) begin 
      x02bai <= 32'b00111111100111101111001010001001;
      x02jyou <= 32'b00111110110001010110000010001110;
    end else if (wbdata[22:12] == 1251) begin 
      x02bai <= 32'b00111111100111101110011000110100;
      x02jyou <= 32'b00111110110001010100000111101110;
    end else if (wbdata[22:12] == 1252) begin 
      x02bai <= 32'b00111111100111101101100111100001;
      x02jyou <= 32'b00111110110001010010001101010110;
    end else if (wbdata[22:12] == 1253) begin 
      x02bai <= 32'b00111111100111101100110110010000;
      x02jyou <= 32'b00111110110001010000010011000110;
    end else if (wbdata[22:12] == 1254) begin 
      x02bai <= 32'b00111111100111101100000101000000;
      x02jyou <= 32'b00111110110001001110011000111010;
    end else if (wbdata[22:12] == 1255) begin 
      x02bai <= 32'b00111111100111101011010011110011;
      x02jyou <= 32'b00111110110001001100011110111000;
    end else if (wbdata[22:12] == 1256) begin 
      x02bai <= 32'b00111111100111101010100010100111;
      x02jyou <= 32'b00111110110001001010100100111010;
    end else if (wbdata[22:12] == 1257) begin 
      x02bai <= 32'b00111111100111101001110001011110;
      x02jyou <= 32'b00111110110001001000101011000111;
    end else if (wbdata[22:12] == 1258) begin 
      x02bai <= 32'b00111111100111101001000000010110;
      x02jyou <= 32'b00111110110001000110110001011001;
    end else if (wbdata[22:12] == 1259) begin 
      x02bai <= 32'b00111111100111101000001111010000;
      x02jyou <= 32'b00111110110001000100110111110001;
    end else if (wbdata[22:12] == 1260) begin 
      x02bai <= 32'b00111111100111100111011110001100;
      x02jyou <= 32'b00111110110001000010111110010001;
    end else if (wbdata[22:12] == 1261) begin 
      x02bai <= 32'b00111111100111100110101101001010;
      x02jyou <= 32'b00111110110001000001000100111001;
    end else if (wbdata[22:12] == 1262) begin 
      x02bai <= 32'b00111111100111100101111100001010;
      x02jyou <= 32'b00111110110000111111001011100111;
    end else if (wbdata[22:12] == 1263) begin 
      x02bai <= 32'b00111111100111100101001011001100;
      x02jyou <= 32'b00111110110000111101010010011101;
    end else if (wbdata[22:12] == 1264) begin 
      x02bai <= 32'b00111111100111100100011010001111;
      x02jyou <= 32'b00111110110000111011011001011000;
    end else if (wbdata[22:12] == 1265) begin 
      x02bai <= 32'b00111111100111100011101001010101;
      x02jyou <= 32'b00111110110000111001100000011100;
    end else if (wbdata[22:12] == 1266) begin 
      x02bai <= 32'b00111111100111100010111000011100;
      x02jyou <= 32'b00111110110000110111100111100110;
    end else if (wbdata[22:12] == 1267) begin 
      x02bai <= 32'b00111111100111100010000111100110;
      x02jyou <= 32'b00111110110000110101101110111001;
    end else if (wbdata[22:12] == 1268) begin 
      x02bai <= 32'b00111111100111100001010110110001;
      x02jyou <= 32'b00111110110000110011110110010001;
    end else if (wbdata[22:12] == 1269) begin 
      x02bai <= 32'b00111111100111100000100101111110;
      x02jyou <= 32'b00111110110000110001111101110000;
    end else if (wbdata[22:12] == 1270) begin 
      x02bai <= 32'b00111111100111011111110101001101;
      x02jyou <= 32'b00111110110000110000000101010110;
    end else if (wbdata[22:12] == 1271) begin 
      x02bai <= 32'b00111111100111011111000100011110;
      x02jyou <= 32'b00111110110000101110001101000100;
    end else if (wbdata[22:12] == 1272) begin 
      x02bai <= 32'b00111111100111011110010011110001;
      x02jyou <= 32'b00111110110000101100010100111001;
    end else if (wbdata[22:12] == 1273) begin 
      x02bai <= 32'b00111111100111011101100011000101;
      x02jyou <= 32'b00111110110000101010011100110010;
    end else if (wbdata[22:12] == 1274) begin 
      x02bai <= 32'b00111111100111011100110010011100;
      x02jyou <= 32'b00111110110000101000100100110110;
    end else if (wbdata[22:12] == 1275) begin 
      x02bai <= 32'b00111111100111011100000001110100;
      x02jyou <= 32'b00111110110000100110101100111110;
    end else if (wbdata[22:12] == 1276) begin 
      x02bai <= 32'b00111111100111011011010001001110;
      x02jyou <= 32'b00111110110000100100110101001101;
    end else if (wbdata[22:12] == 1277) begin 
      x02bai <= 32'b00111111100111011010100000101010;
      x02jyou <= 32'b00111110110000100010111101100100;
    end else if (wbdata[22:12] == 1278) begin 
      x02bai <= 32'b00111111100111011001110000001000;
      x02jyou <= 32'b00111110110000100001000110000010;
    end else if (wbdata[22:12] == 1279) begin 
      x02bai <= 32'b00111111100111011000111111101000;
      x02jyou <= 32'b00111110110000011111001110100111;
    end else if (wbdata[22:12] == 1280) begin 
      x02bai <= 32'b00111111100111011000001111001010;
      x02jyou <= 32'b00111110110000011101010111010011;
    end else if (wbdata[22:12] == 1281) begin 
      x02bai <= 32'b00111111100111010111011110101110;
      x02jyou <= 32'b00111110110000011011100000000111;
    end else if (wbdata[22:12] == 1282) begin 
      x02bai <= 32'b00111111100111010110101110010011;
      x02jyou <= 32'b00111110110000011001101000111111;
    end else if (wbdata[22:12] == 1283) begin 
      x02bai <= 32'b00111111100111010101111101111010;
      x02jyou <= 32'b00111110110000010111110001111110;
    end else if (wbdata[22:12] == 1284) begin 
      x02bai <= 32'b00111111100111010101001101100011;
      x02jyou <= 32'b00111110110000010101111011000101;
    end else if (wbdata[22:12] == 1285) begin 
      x02bai <= 32'b00111111100111010100011101001110;
      x02jyou <= 32'b00111110110000010100000100010011;
    end else if (wbdata[22:12] == 1286) begin 
      x02bai <= 32'b00111111100111010011101100111011;
      x02jyou <= 32'b00111110110000010010001101101000;
    end else if (wbdata[22:12] == 1287) begin 
      x02bai <= 32'b00111111100111010010111100101010;
      x02jyou <= 32'b00111110110000010000010111000100;
    end else if (wbdata[22:12] == 1288) begin 
      x02bai <= 32'b00111111100111010010001100011011;
      x02jyou <= 32'b00111110110000001110100000101000;
    end else if (wbdata[22:12] == 1289) begin 
      x02bai <= 32'b00111111100111010001011100001101;
      x02jyou <= 32'b00111110110000001100101010010000;
    end else if (wbdata[22:12] == 1290) begin 
      x02bai <= 32'b00111111100111010000101100000001;
      x02jyou <= 32'b00111110110000001010110011111111;
    end else if (wbdata[22:12] == 1291) begin 
      x02bai <= 32'b00111111100111001111111011110111;
      x02jyou <= 32'b00111110110000001000111101110110;
    end else if (wbdata[22:12] == 1292) begin 
      x02bai <= 32'b00111111100111001111001011101111;
      x02jyou <= 32'b00111110110000000111000111110100;
    end else if (wbdata[22:12] == 1293) begin 
      x02bai <= 32'b00111111100111001110011011101001;
      x02jyou <= 32'b00111110110000000101010001111000;
    end else if (wbdata[22:12] == 1294) begin 
      x02bai <= 32'b00111111100111001101101011100101;
      x02jyou <= 32'b00111110110000000011011100000101;
    end else if (wbdata[22:12] == 1295) begin 
      x02bai <= 32'b00111111100111001100111011100010;
      x02jyou <= 32'b00111110110000000001100110010101;
    end else if (wbdata[22:12] == 1296) begin 
      x02bai <= 32'b00111111100111001100001011100001;
      x02jyou <= 32'b00111110101111111111110000101101;
    end else if (wbdata[22:12] == 1297) begin 
      x02bai <= 32'b00111111100111001011011011100011;
      x02jyou <= 32'b00111110101111111101111011001111;
    end else if (wbdata[22:12] == 1298) begin 
      x02bai <= 32'b00111111100111001010101011100110;
      x02jyou <= 32'b00111110101111111100000101110101;
    end else if (wbdata[22:12] == 1299) begin 
      x02bai <= 32'b00111111100111001001111011101010;
      x02jyou <= 32'b00111110101111111010010000100000;
    end else if (wbdata[22:12] == 1300) begin 
      x02bai <= 32'b00111111100111001001001011110001;
      x02jyou <= 32'b00111110101111111000011011010100;
    end else if (wbdata[22:12] == 1301) begin 
      x02bai <= 32'b00111111100111001000011011111010;
      x02jyou <= 32'b00111110101111110110100110010000;
    end else if (wbdata[22:12] == 1302) begin 
      x02bai <= 32'b00111111100111000111101100000100;
      x02jyou <= 32'b00111110101111110100110001010000;
    end else if (wbdata[22:12] == 1303) begin 
      x02bai <= 32'b00111111100111000110111100010000;
      x02jyou <= 32'b00111110101111110010111100010111;
    end else if (wbdata[22:12] == 1304) begin 
      x02bai <= 32'b00111111100111000110001100011110;
      x02jyou <= 32'b00111110101111110001000111100110;
    end else if (wbdata[22:12] == 1305) begin 
      x02bai <= 32'b00111111100111000101011100101110;
      x02jyou <= 32'b00111110101111101111010010111100;
    end else if (wbdata[22:12] == 1306) begin 
      x02bai <= 32'b00111111100111000100101100111111;
      x02jyou <= 32'b00111110101111101101011110010110;
    end else if (wbdata[22:12] == 1307) begin 
      x02bai <= 32'b00111111100111000011111101010011;
      x02jyou <= 32'b00111110101111101011101001111010;
    end else if (wbdata[22:12] == 1308) begin 
      x02bai <= 32'b00111111100111000011001101101000;
      x02jyou <= 32'b00111110101111101001110101100010;
    end else if (wbdata[22:12] == 1309) begin 
      x02bai <= 32'b00111111100111000010011101111111;
      x02jyou <= 32'b00111110101111101000000001010010;
    end else if (wbdata[22:12] == 1310) begin 
      x02bai <= 32'b00111111100111000001101110011000;
      x02jyou <= 32'b00111110101111100110001101001000;
    end else if (wbdata[22:12] == 1311) begin 
      x02bai <= 32'b00111111100111000000111110110011;
      x02jyou <= 32'b00111110101111100100011001000110;
    end else if (wbdata[22:12] == 1312) begin 
      x02bai <= 32'b00111111100111000000001111001111;
      x02jyou <= 32'b00111110101111100010100101001001;
    end else if (wbdata[22:12] == 1313) begin 
      x02bai <= 32'b00111111100110111111011111101110;
      x02jyou <= 32'b00111110101111100000110001010101;
    end else if (wbdata[22:12] == 1314) begin 
      x02bai <= 32'b00111111100110111110110000001110;
      x02jyou <= 32'b00111110101111011110111101100101;
    end else if (wbdata[22:12] == 1315) begin 
      x02bai <= 32'b00111111100110111110000000110000;
      x02jyou <= 32'b00111110101111011101001001111101;
    end else if (wbdata[22:12] == 1316) begin 
      x02bai <= 32'b00111111100110111101010001010011;
      x02jyou <= 32'b00111110101111011011010110011001;
    end else if (wbdata[22:12] == 1317) begin 
      x02bai <= 32'b00111111100110111100100001111001;
      x02jyou <= 32'b00111110101111011001100010111111;
    end else if (wbdata[22:12] == 1318) begin 
      x02bai <= 32'b00111111100110111011110010100000;
      x02jyou <= 32'b00111110101111010111101111101001;
    end else if (wbdata[22:12] == 1319) begin 
      x02bai <= 32'b00111111100110111011000011001010;
      x02jyou <= 32'b00111110101111010101111100011101;
    end else if (wbdata[22:12] == 1320) begin 
      x02bai <= 32'b00111111100110111010010011110100;
      x02jyou <= 32'b00111110101111010100001001010100;
    end else if (wbdata[22:12] == 1321) begin 
      x02bai <= 32'b00111111100110111001100100100001;
      x02jyou <= 32'b00111110101111010010010110010011;
    end else if (wbdata[22:12] == 1322) begin 
      x02bai <= 32'b00111111100110111000110101010000;
      x02jyou <= 32'b00111110101111010000100011011010;
    end else if (wbdata[22:12] == 1323) begin 
      x02bai <= 32'b00111111100110111000000110000000;
      x02jyou <= 32'b00111110101111001110110000100101;
    end else if (wbdata[22:12] == 1324) begin 
      x02bai <= 32'b00111111100110110111010110110010;
      x02jyou <= 32'b00111110101111001100111101110111;
    end else if (wbdata[22:12] == 1325) begin 
      x02bai <= 32'b00111111100110110110100111100110;
      x02jyou <= 32'b00111110101111001011001011010001;
    end else if (wbdata[22:12] == 1326) begin 
      x02bai <= 32'b00111111100110110101111000011100;
      x02jyou <= 32'b00111110101111001001011000110001;
    end else if (wbdata[22:12] == 1327) begin 
      x02bai <= 32'b00111111100110110101001001010011;
      x02jyou <= 32'b00111110101111000111100110010110;
    end else if (wbdata[22:12] == 1328) begin 
      x02bai <= 32'b00111111100110110100011010001101;
      x02jyou <= 32'b00111110101111000101110100000100;
    end else if (wbdata[22:12] == 1329) begin 
      x02bai <= 32'b00111111100110110011101011001000;
      x02jyou <= 32'b00111110101111000100000001110111;
    end else if (wbdata[22:12] == 1330) begin 
      x02bai <= 32'b00111111100110110010111100000101;
      x02jyou <= 32'b00111110101111000010001111110001;
    end else if (wbdata[22:12] == 1331) begin 
      x02bai <= 32'b00111111100110110010001101000011;
      x02jyou <= 32'b00111110101111000000011101110000;
    end else if (wbdata[22:12] == 1332) begin 
      x02bai <= 32'b00111111100110110001011110000100;
      x02jyou <= 32'b00111110101110111110101011111000;
    end else if (wbdata[22:12] == 1333) begin 
      x02bai <= 32'b00111111100110110000101111000110;
      x02jyou <= 32'b00111110101110111100111010000101;
    end else if (wbdata[22:12] == 1334) begin 
      x02bai <= 32'b00111111100110110000000000001010;
      x02jyou <= 32'b00111110101110111011001000011000;
    end else if (wbdata[22:12] == 1335) begin 
      x02bai <= 32'b00111111100110101111010001010000;
      x02jyou <= 32'b00111110101110111001010110110011;
    end else if (wbdata[22:12] == 1336) begin 
      x02bai <= 32'b00111111100110101110100010010111;
      x02jyou <= 32'b00111110101110110111100101010010;
    end else if (wbdata[22:12] == 1337) begin 
      x02bai <= 32'b00111111100110101101110011100001;
      x02jyou <= 32'b00111110101110110101110011111011;
    end else if (wbdata[22:12] == 1338) begin 
      x02bai <= 32'b00111111100110101101000100101100;
      x02jyou <= 32'b00111110101110110100000010101000;
    end else if (wbdata[22:12] == 1339) begin 
      x02bai <= 32'b00111111100110101100010101111000;
      x02jyou <= 32'b00111110101110110010010001011001;
    end else if (wbdata[22:12] == 1340) begin 
      x02bai <= 32'b00111111100110101011100111000111;
      x02jyou <= 32'b00111110101110110000100000010100;
    end else if (wbdata[22:12] == 1341) begin 
      x02bai <= 32'b00111111100110101010111000010111;
      x02jyou <= 32'b00111110101110101110101111010100;
    end else if (wbdata[22:12] == 1342) begin 
      x02bai <= 32'b00111111100110101010001001101010;
      x02jyou <= 32'b00111110101110101100111110011101;
    end else if (wbdata[22:12] == 1343) begin 
      x02bai <= 32'b00111111100110101001011010111101;
      x02jyou <= 32'b00111110101110101011001101101000;
    end else if (wbdata[22:12] == 1344) begin 
      x02bai <= 32'b00111111100110101000101100010011;
      x02jyou <= 32'b00111110101110101001011100111101;
    end else if (wbdata[22:12] == 1345) begin 
      x02bai <= 32'b00111111100110100111111101101011;
      x02jyou <= 32'b00111110101110100111101100011000;
    end else if (wbdata[22:12] == 1346) begin 
      x02bai <= 32'b00111111100110100111001111000100;
      x02jyou <= 32'b00111110101110100101111011111000;
    end else if (wbdata[22:12] == 1347) begin 
      x02bai <= 32'b00111111100110100110100000011111;
      x02jyou <= 32'b00111110101110100100001011011111;
    end else if (wbdata[22:12] == 1348) begin 
      x02bai <= 32'b00111111100110100101110001111011;
      x02jyou <= 32'b00111110101110100010011011001011;
    end else if (wbdata[22:12] == 1349) begin 
      x02bai <= 32'b00111111100110100101000011011010;
      x02jyou <= 32'b00111110101110100000101011000000;
    end else if (wbdata[22:12] == 1350) begin 
      x02bai <= 32'b00111111100110100100010100111010;
      x02jyou <= 32'b00111110101110011110111010111001;
    end else if (wbdata[22:12] == 1351) begin 
      x02bai <= 32'b00111111100110100011100110011100;
      x02jyou <= 32'b00111110101110011101001010111001;
    end else if (wbdata[22:12] == 1352) begin 
      x02bai <= 32'b00111111100110100010111000000000;
      x02jyou <= 32'b00111110101110011011011011000001;
    end else if (wbdata[22:12] == 1353) begin 
      x02bai <= 32'b00111111100110100010001001100101;
      x02jyou <= 32'b00111110101110011001101011001100;
    end else if (wbdata[22:12] == 1354) begin 
      x02bai <= 32'b00111111100110100001011011001100;
      x02jyou <= 32'b00111110101110010111111011011111;
    end else if (wbdata[22:12] == 1355) begin 
      x02bai <= 32'b00111111100110100000101100110101;
      x02jyou <= 32'b00111110101110010110001011111001;
    end else if (wbdata[22:12] == 1356) begin 
      x02bai <= 32'b00111111100110011111111110100000;
      x02jyou <= 32'b00111110101110010100011100011001;
    end else if (wbdata[22:12] == 1357) begin 
      x02bai <= 32'b00111111100110011111010000001100;
      x02jyou <= 32'b00111110101110010010101100111110;
    end else if (wbdata[22:12] == 1358) begin 
      x02bai <= 32'b00111111100110011110100001111011;
      x02jyou <= 32'b00111110101110010000111101101100;
    end else if (wbdata[22:12] == 1359) begin 
      x02bai <= 32'b00111111100110011101110011101010;
      x02jyou <= 32'b00111110101110001111001110011101;
    end else if (wbdata[22:12] == 1360) begin 
      x02bai <= 32'b00111111100110011101000101011100;
      x02jyou <= 32'b00111110101110001101011111010110;
    end else if (wbdata[22:12] == 1361) begin 
      x02bai <= 32'b00111111100110011100010111001111;
      x02jyou <= 32'b00111110101110001011110000010101;
    end else if (wbdata[22:12] == 1362) begin 
      x02bai <= 32'b00111111100110011011101001000101;
      x02jyou <= 32'b00111110101110001010000001011100;
    end else if (wbdata[22:12] == 1363) begin 
      x02bai <= 32'b00111111100110011010111010111011;
      x02jyou <= 32'b00111110101110001000010010100110;
    end else if (wbdata[22:12] == 1364) begin 
      x02bai <= 32'b00111111100110011010001100110100;
      x02jyou <= 32'b00111110101110000110100011111000;
    end else if (wbdata[22:12] == 1365) begin 
      x02bai <= 32'b00111111100110011001011110101110;
      x02jyou <= 32'b00111110101110000100110101010000;
    end else if (wbdata[22:12] == 1366) begin 
      x02bai <= 32'b00111111100110011000110000101010;
      x02jyou <= 32'b00111110101110000011000110101110;
    end else if (wbdata[22:12] == 1367) begin 
      x02bai <= 32'b00111111100110011000000010101000;
      x02jyou <= 32'b00111110101110000001011000010011;
    end else if (wbdata[22:12] == 1368) begin 
      x02bai <= 32'b00111111100110010111010100101000;
      x02jyou <= 32'b00111110101101111111101001111111;
    end else if (wbdata[22:12] == 1369) begin 
      x02bai <= 32'b00111111100110010110100110101001;
      x02jyou <= 32'b00111110101101111101111011101111;
    end else if (wbdata[22:12] == 1370) begin 
      x02bai <= 32'b00111111100110010101111000101100;
      x02jyou <= 32'b00111110101101111100001101100110;
    end else if (wbdata[22:12] == 1371) begin 
      x02bai <= 32'b00111111100110010101001010110000;
      x02jyou <= 32'b00111110101101111010011111100010;
    end else if (wbdata[22:12] == 1372) begin 
      x02bai <= 32'b00111111100110010100011100110111;
      x02jyou <= 32'b00111110101101111000110001100111;
    end else if (wbdata[22:12] == 1373) begin 
      x02bai <= 32'b00111111100110010011101110111111;
      x02jyou <= 32'b00111110101101110111000011110000;
    end else if (wbdata[22:12] == 1374) begin 
      x02bai <= 32'b00111111100110010011000001001001;
      x02jyou <= 32'b00111110101101110101010110000001;
    end else if (wbdata[22:12] == 1375) begin 
      x02bai <= 32'b00111111100110010010010011010100;
      x02jyou <= 32'b00111110101101110011101000010101;
    end else if (wbdata[22:12] == 1376) begin 
      x02bai <= 32'b00111111100110010001100101100001;
      x02jyou <= 32'b00111110101101110001111010110001;
    end else if (wbdata[22:12] == 1377) begin 
      x02bai <= 32'b00111111100110010000110111110000;
      x02jyou <= 32'b00111110101101110000001101010011;
    end else if (wbdata[22:12] == 1378) begin 
      x02bai <= 32'b00111111100110010000001010000001;
      x02jyou <= 32'b00111110101101101110011111111100;
    end else if (wbdata[22:12] == 1379) begin 
      x02bai <= 32'b00111111100110001111011100010011;
      x02jyou <= 32'b00111110101101101100110010101010;
    end else if (wbdata[22:12] == 1380) begin 
      x02bai <= 32'b00111111100110001110101110100111;
      x02jyou <= 32'b00111110101101101011000101011110;
    end else if (wbdata[22:12] == 1381) begin 
      x02bai <= 32'b00111111100110001110000000111101;
      x02jyou <= 32'b00111110101101101001011000011010;
    end else if (wbdata[22:12] == 1382) begin 
      x02bai <= 32'b00111111100110001101010011010101;
      x02jyou <= 32'b00111110101101100111101011011100;
    end else if (wbdata[22:12] == 1383) begin 
      x02bai <= 32'b00111111100110001100100101101110;
      x02jyou <= 32'b00111110101101100101111110100010;
    end else if (wbdata[22:12] == 1384) begin 
      x02bai <= 32'b00111111100110001011111000001001;
      x02jyou <= 32'b00111110101101100100010001110000;
    end else if (wbdata[22:12] == 1385) begin 
      x02bai <= 32'b00111111100110001011001010100101;
      x02jyou <= 32'b00111110101101100010100101000001;
    end else if (wbdata[22:12] == 1386) begin 
      x02bai <= 32'b00111111100110001010011101000011;
      x02jyou <= 32'b00111110101101100000111000011010;
    end else if (wbdata[22:12] == 1387) begin 
      x02bai <= 32'b00111111100110001001101111100011;
      x02jyou <= 32'b00111110101101011111001011111001;
    end else if (wbdata[22:12] == 1388) begin 
      x02bai <= 32'b00111111100110001001000010000101;
      x02jyou <= 32'b00111110101101011101011111011111;
    end else if (wbdata[22:12] == 1389) begin 
      x02bai <= 32'b00111111100110001000010100101000;
      x02jyou <= 32'b00111110101101011011110011001010;
    end else if (wbdata[22:12] == 1390) begin 
      x02bai <= 32'b00111111100110000111100111001110;
      x02jyou <= 32'b00111110101101011010000110111101;
    end else if (wbdata[22:12] == 1391) begin 
      x02bai <= 32'b00111111100110000110111001110100;
      x02jyou <= 32'b00111110101101011000011010110011;
    end else if (wbdata[22:12] == 1392) begin 
      x02bai <= 32'b00111111100110000110001100011101;
      x02jyou <= 32'b00111110101101010110101110110010;
    end else if (wbdata[22:12] == 1393) begin 
      x02bai <= 32'b00111111100110000101011111000111;
      x02jyou <= 32'b00111110101101010101000010110101;
    end else if (wbdata[22:12] == 1394) begin 
      x02bai <= 32'b00111111100110000100110001110011;
      x02jyou <= 32'b00111110101101010011010110111111;
    end else if (wbdata[22:12] == 1395) begin 
      x02bai <= 32'b00111111100110000100000100100000;
      x02jyou <= 32'b00111110101101010001101011001101;
    end else if (wbdata[22:12] == 1396) begin 
      x02bai <= 32'b00111111100110000011010111001111;
      x02jyou <= 32'b00111110101101001111111111100010;
    end else if (wbdata[22:12] == 1397) begin 
      x02bai <= 32'b00111111100110000010101010000000;
      x02jyou <= 32'b00111110101101001110010011111110;
    end else if (wbdata[22:12] == 1398) begin 
      x02bai <= 32'b00111111100110000001111100110011;
      x02jyou <= 32'b00111110101101001100101000100001;
    end else if (wbdata[22:12] == 1399) begin 
      x02bai <= 32'b00111111100110000001001111100111;
      x02jyou <= 32'b00111110101101001010111101001000;
    end else if (wbdata[22:12] == 1400) begin 
      x02bai <= 32'b00111111100110000000100010011101;
      x02jyou <= 32'b00111110101101001001010001110101;
    end else if (wbdata[22:12] == 1401) begin 
      x02bai <= 32'b00111111100101111111110101010100;
      x02jyou <= 32'b00111110101101000111100110101000;
    end else if (wbdata[22:12] == 1402) begin 
      x02bai <= 32'b00111111100101111111001000001101;
      x02jyou <= 32'b00111110101101000101111011100000;
    end else if (wbdata[22:12] == 1403) begin 
      x02bai <= 32'b00111111100101111110011011001000;
      x02jyou <= 32'b00111110101101000100010000100000;
    end else if (wbdata[22:12] == 1404) begin 
      x02bai <= 32'b00111111100101111101101110000101;
      x02jyou <= 32'b00111110101101000010100101100110;
    end else if (wbdata[22:12] == 1405) begin 
      x02bai <= 32'b00111111100101111101000001000011;
      x02jyou <= 32'b00111110101101000000111010110001;
    end else if (wbdata[22:12] == 1406) begin 
      x02bai <= 32'b00111111100101111100010100000011;
      x02jyou <= 32'b00111110101100111111010000000010;
    end else if (wbdata[22:12] == 1407) begin 
      x02bai <= 32'b00111111100101111011100111000101;
      x02jyou <= 32'b00111110101100111101100101011010;
    end else if (wbdata[22:12] == 1408) begin 
      x02bai <= 32'b00111111100101111010111010001000;
      x02jyou <= 32'b00111110101100111011111010110111;
    end else if (wbdata[22:12] == 1409) begin 
      x02bai <= 32'b00111111100101111010001101001101;
      x02jyou <= 32'b00111110101100111010010000011010;
    end else if (wbdata[22:12] == 1410) begin 
      x02bai <= 32'b00111111100101111001100000010011;
      x02jyou <= 32'b00111110101100111000100110000010;
    end else if (wbdata[22:12] == 1411) begin 
      x02bai <= 32'b00111111100101111000110011011100;
      x02jyou <= 32'b00111110101100110110111011110010;
    end else if (wbdata[22:12] == 1412) begin 
      x02bai <= 32'b00111111100101111000000110100110;
      x02jyou <= 32'b00111110101100110101010001100111;
    end else if (wbdata[22:12] == 1413) begin 
      x02bai <= 32'b00111111100101110111011001110001;
      x02jyou <= 32'b00111110101100110011100111100000;
    end else if (wbdata[22:12] == 1414) begin 
      x02bai <= 32'b00111111100101110110101100111110;
      x02jyou <= 32'b00111110101100110001111101100000;
    end else if (wbdata[22:12] == 1415) begin 
      x02bai <= 32'b00111111100101110110000000001101;
      x02jyou <= 32'b00111110101100110000010011100111;
    end else if (wbdata[22:12] == 1416) begin 
      x02bai <= 32'b00111111100101110101010011011110;
      x02jyou <= 32'b00111110101100101110101001110100;
    end else if (wbdata[22:12] == 1417) begin 
      x02bai <= 32'b00111111100101110100100110110000;
      x02jyou <= 32'b00111110101100101101000000000110;
    end else if (wbdata[22:12] == 1418) begin 
      x02bai <= 32'b00111111100101110011111010000100;
      x02jyou <= 32'b00111110101100101011010110011110;
    end else if (wbdata[22:12] == 1419) begin 
      x02bai <= 32'b00111111100101110011001101011001;
      x02jyou <= 32'b00111110101100101001101100111011;
    end else if (wbdata[22:12] == 1420) begin 
      x02bai <= 32'b00111111100101110010100000110000;
      x02jyou <= 32'b00111110101100101000000011011110;
    end else if (wbdata[22:12] == 1421) begin 
      x02bai <= 32'b00111111100101110001110100001001;
      x02jyou <= 32'b00111110101100100110011010001000;
    end else if (wbdata[22:12] == 1422) begin 
      x02bai <= 32'b00111111100101110001000111100100;
      x02jyou <= 32'b00111110101100100100110000111000;
    end else if (wbdata[22:12] == 1423) begin 
      x02bai <= 32'b00111111100101110000011011000000;
      x02jyou <= 32'b00111110101100100011000111101101;
    end else if (wbdata[22:12] == 1424) begin 
      x02bai <= 32'b00111111100101101111101110011101;
      x02jyou <= 32'b00111110101100100001011110100111;
    end else if (wbdata[22:12] == 1425) begin 
      x02bai <= 32'b00111111100101101111000001111101;
      x02jyou <= 32'b00111110101100011111110101101001;
    end else if (wbdata[22:12] == 1426) begin 
      x02bai <= 32'b00111111100101101110010101011110;
      x02jyou <= 32'b00111110101100011110001100101111;
    end else if (wbdata[22:12] == 1427) begin 
      x02bai <= 32'b00111111100101101101101001000000;
      x02jyou <= 32'b00111110101100011100100011111010;
    end else if (wbdata[22:12] == 1428) begin 
      x02bai <= 32'b00111111100101101100111100100100;
      x02jyou <= 32'b00111110101100011010111011001100;
    end else if (wbdata[22:12] == 1429) begin 
      x02bai <= 32'b00111111100101101100010000001010;
      x02jyou <= 32'b00111110101100011001010010100100;
    end else if (wbdata[22:12] == 1430) begin 
      x02bai <= 32'b00111111100101101011100011110010;
      x02jyou <= 32'b00111110101100010111101010000010;
    end else if (wbdata[22:12] == 1431) begin 
      x02bai <= 32'b00111111100101101010110111011011;
      x02jyou <= 32'b00111110101100010110000001100101;
    end else if (wbdata[22:12] == 1432) begin 
      x02bai <= 32'b00111111100101101010001011000110;
      x02jyou <= 32'b00111110101100010100011001001111;
    end else if (wbdata[22:12] == 1433) begin 
      x02bai <= 32'b00111111100101101001011110110010;
      x02jyou <= 32'b00111110101100010010110000111101;
    end else if (wbdata[22:12] == 1434) begin 
      x02bai <= 32'b00111111100101101000110010100000;
      x02jyou <= 32'b00111110101100010001001000110001;
    end else if (wbdata[22:12] == 1435) begin 
      x02bai <= 32'b00111111100101101000000110010000;
      x02jyou <= 32'b00111110101100001111100000101101;
    end else if (wbdata[22:12] == 1436) begin 
      x02bai <= 32'b00111111100101100111011010000001;
      x02jyou <= 32'b00111110101100001101111000101100;
    end else if (wbdata[22:12] == 1437) begin 
      x02bai <= 32'b00111111100101100110101101110100;
      x02jyou <= 32'b00111110101100001100010000110010;
    end else if (wbdata[22:12] == 1438) begin 
      x02bai <= 32'b00111111100101100110000001101001;
      x02jyou <= 32'b00111110101100001010101000111111;
    end else if (wbdata[22:12] == 1439) begin 
      x02bai <= 32'b00111111100101100101010101011111;
      x02jyou <= 32'b00111110101100001001000001010000;
    end else if (wbdata[22:12] == 1440) begin 
      x02bai <= 32'b00111111100101100100101001010111;
      x02jyou <= 32'b00111110101100000111011001100111;
    end else if (wbdata[22:12] == 1441) begin 
      x02bai <= 32'b00111111100101100011111101010000;
      x02jyou <= 32'b00111110101100000101110010000011;
    end else if (wbdata[22:12] == 1442) begin 
      x02bai <= 32'b00111111100101100011010001001011;
      x02jyou <= 32'b00111110101100000100001010100101;
    end else if (wbdata[22:12] == 1443) begin 
      x02bai <= 32'b00111111100101100010100101001000;
      x02jyou <= 32'b00111110101100000010100011001110;
    end else if (wbdata[22:12] == 1444) begin 
      x02bai <= 32'b00111111100101100001111001000110;
      x02jyou <= 32'b00111110101100000000111011111011;
    end else if (wbdata[22:12] == 1445) begin 
      x02bai <= 32'b00111111100101100001001101000110;
      x02jyou <= 32'b00111110101011111111010100101111;
    end else if (wbdata[22:12] == 1446) begin 
      x02bai <= 32'b00111111100101100000100001000111;
      x02jyou <= 32'b00111110101011111101101101100111;
    end else if (wbdata[22:12] == 1447) begin 
      x02bai <= 32'b00111111100101011111110101001011;
      x02jyou <= 32'b00111110101011111100000110101000;
    end else if (wbdata[22:12] == 1448) begin 
      x02bai <= 32'b00111111100101011111001001001111;
      x02jyou <= 32'b00111110101011111010011111101011;
    end else if (wbdata[22:12] == 1449) begin 
      x02bai <= 32'b00111111100101011110011101010110;
      x02jyou <= 32'b00111110101011111000111000110110;
    end else if (wbdata[22:12] == 1450) begin 
      x02bai <= 32'b00111111100101011101110001011101;
      x02jyou <= 32'b00111110101011110111010010000100;
    end else if (wbdata[22:12] == 1451) begin 
      x02bai <= 32'b00111111100101011101000101100111;
      x02jyou <= 32'b00111110101011110101101011011010;
    end else if (wbdata[22:12] == 1452) begin 
      x02bai <= 32'b00111111100101011100011001110010;
      x02jyou <= 32'b00111110101011110100000100110101;
    end else if (wbdata[22:12] == 1453) begin 
      x02bai <= 32'b00111111100101011011101101111111;
      x02jyou <= 32'b00111110101011110010011110010110;
    end else if (wbdata[22:12] == 1454) begin 
      x02bai <= 32'b00111111100101011011000010001101;
      x02jyou <= 32'b00111110101011110000110111111100;
    end else if (wbdata[22:12] == 1455) begin 
      x02bai <= 32'b00111111100101011010010110011101;
      x02jyou <= 32'b00111110101011101111010001101000;
    end else if (wbdata[22:12] == 1456) begin 
      x02bai <= 32'b00111111100101011001101010101111;
      x02jyou <= 32'b00111110101011101101101011011010;
    end else if (wbdata[22:12] == 1457) begin 
      x02bai <= 32'b00111111100101011000111111000010;
      x02jyou <= 32'b00111110101011101100000101010001;
    end else if (wbdata[22:12] == 1458) begin 
      x02bai <= 32'b00111111100101011000010011010110;
      x02jyou <= 32'b00111110101011101010011111001100;
    end else if (wbdata[22:12] == 1459) begin 
      x02bai <= 32'b00111111100101010111100111101101;
      x02jyou <= 32'b00111110101011101000111001010000;
    end else if (wbdata[22:12] == 1460) begin 
      x02bai <= 32'b00111111100101010110111100000101;
      x02jyou <= 32'b00111110101011100111010011011000;
    end else if (wbdata[22:12] == 1461) begin 
      x02bai <= 32'b00111111100101010110010000011110;
      x02jyou <= 32'b00111110101011100101101101100100;
    end else if (wbdata[22:12] == 1462) begin 
      x02bai <= 32'b00111111100101010101100100111001;
      x02jyou <= 32'b00111110101011100100000111110111;
    end else if (wbdata[22:12] == 1463) begin 
      x02bai <= 32'b00111111100101010100111001010110;
      x02jyou <= 32'b00111110101011100010100010010000;
    end else if (wbdata[22:12] == 1464) begin 
      x02bai <= 32'b00111111100101010100001101110100;
      x02jyou <= 32'b00111110101011100000111100101110;
    end else if (wbdata[22:12] == 1465) begin 
      x02bai <= 32'b00111111100101010011100010010100;
      x02jyou <= 32'b00111110101011011111010111010010;
    end else if (wbdata[22:12] == 1466) begin 
      x02bai <= 32'b00111111100101010010110110110101;
      x02jyou <= 32'b00111110101011011101110001111010;
    end else if (wbdata[22:12] == 1467) begin 
      x02bai <= 32'b00111111100101010010001011011000;
      x02jyou <= 32'b00111110101011011100001100101000;
    end else if (wbdata[22:12] == 1468) begin 
      x02bai <= 32'b00111111100101010001011111111101;
      x02jyou <= 32'b00111110101011011010100111011110;
    end else if (wbdata[22:12] == 1469) begin 
      x02bai <= 32'b00111111100101010000110100100011;
      x02jyou <= 32'b00111110101011011001000010010111;
    end else if (wbdata[22:12] == 1470) begin 
      x02bai <= 32'b00111111100101010000001001001011;
      x02jyou <= 32'b00111110101011010111011101010111;
    end else if (wbdata[22:12] == 1471) begin 
      x02bai <= 32'b00111111100101001111011101110100;
      x02jyou <= 32'b00111110101011010101111000011011;
    end else if (wbdata[22:12] == 1472) begin 
      x02bai <= 32'b00111111100101001110110010011111;
      x02jyou <= 32'b00111110101011010100010011100101;
    end else if (wbdata[22:12] == 1473) begin 
      x02bai <= 32'b00111111100101001110000111001100;
      x02jyou <= 32'b00111110101011010010101110110110;
    end else if (wbdata[22:12] == 1474) begin 
      x02bai <= 32'b00111111100101001101011011111010;
      x02jyou <= 32'b00111110101011010001001010001011;
    end else if (wbdata[22:12] == 1475) begin 
      x02bai <= 32'b00111111100101001100110000101001;
      x02jyou <= 32'b00111110101011001111100101100100;
    end else if (wbdata[22:12] == 1476) begin 
      x02bai <= 32'b00111111100101001100000101011011;
      x02jyou <= 32'b00111110101011001110000001000111;
    end else if (wbdata[22:12] == 1477) begin 
      x02bai <= 32'b00111111100101001011011010001101;
      x02jyou <= 32'b00111110101011001100011100101010;
    end else if (wbdata[22:12] == 1478) begin 
      x02bai <= 32'b00111111100101001010101111000010;
      x02jyou <= 32'b00111110101011001010111000010111;
    end else if (wbdata[22:12] == 1479) begin 
      x02bai <= 32'b00111111100101001010000011111000;
      x02jyou <= 32'b00111110101011001001010100001000;
    end else if (wbdata[22:12] == 1480) begin 
      x02bai <= 32'b00111111100101001001011000101111;
      x02jyou <= 32'b00111110101011000111101111111101;
    end else if (wbdata[22:12] == 1481) begin 
      x02bai <= 32'b00111111100101001000101101101000;
      x02jyou <= 32'b00111110101011000110001011111000;
    end else if (wbdata[22:12] == 1482) begin 
      x02bai <= 32'b00111111100101001000000010100011;
      x02jyou <= 32'b00111110101011000100100111111010;
    end else if (wbdata[22:12] == 1483) begin 
      x02bai <= 32'b00111111100101000111010111011111;
      x02jyou <= 32'b00111110101011000011000100000000;
    end else if (wbdata[22:12] == 1484) begin 
      x02bai <= 32'b00111111100101000110101100011100;
      x02jyou <= 32'b00111110101011000001100000001010;
    end else if (wbdata[22:12] == 1485) begin 
      x02bai <= 32'b00111111100101000110000001011100;
      x02jyou <= 32'b00111110101010111111111100011101;
    end else if (wbdata[22:12] == 1486) begin 
      x02bai <= 32'b00111111100101000101010110011101;
      x02jyou <= 32'b00111110101010111110011000110100;
    end else if (wbdata[22:12] == 1487) begin 
      x02bai <= 32'b00111111100101000100101011011111;
      x02jyou <= 32'b00111110101010111100110101001111;
    end else if (wbdata[22:12] == 1488) begin 
      x02bai <= 32'b00111111100101000100000000100011;
      x02jyou <= 32'b00111110101010111011010001110001;
    end else if (wbdata[22:12] == 1489) begin 
      x02bai <= 32'b00111111100101000011010101101000;
      x02jyou <= 32'b00111110101010111001101110010111;
    end else if (wbdata[22:12] == 1490) begin 
      x02bai <= 32'b00111111100101000010101010101111;
      x02jyou <= 32'b00111110101010111000001011000011;
    end else if (wbdata[22:12] == 1491) begin 
      x02bai <= 32'b00111111100101000001111111111000;
      x02jyou <= 32'b00111110101010110110100111110101;
    end else if (wbdata[22:12] == 1492) begin 
      x02bai <= 32'b00111111100101000001010101000010;
      x02jyou <= 32'b00111110101010110101000100101100;
    end else if (wbdata[22:12] == 1493) begin 
      x02bai <= 32'b00111111100101000000101010001110;
      x02jyou <= 32'b00111110101010110011100001101001;
    end else if (wbdata[22:12] == 1494) begin 
      x02bai <= 32'b00111111100100111111111111011011;
      x02jyou <= 32'b00111110101010110001111110101010;
    end else if (wbdata[22:12] == 1495) begin 
      x02bai <= 32'b00111111100100111111010100101010;
      x02jyou <= 32'b00111110101010110000011011110010;
    end else if (wbdata[22:12] == 1496) begin 
      x02bai <= 32'b00111111100100111110101001111010;
      x02jyou <= 32'b00111110101010101110111000111110;
    end else if (wbdata[22:12] == 1497) begin 
      x02bai <= 32'b00111111100100111101111111001100;
      x02jyou <= 32'b00111110101010101101010110010000;
    end else if (wbdata[22:12] == 1498) begin 
      x02bai <= 32'b00111111100100111101010100100000;
      x02jyou <= 32'b00111110101010101011110011101000;
    end else if (wbdata[22:12] == 1499) begin 
      x02bai <= 32'b00111111100100111100101001110101;
      x02jyou <= 32'b00111110101010101010010001000101;
    end else if (wbdata[22:12] == 1500) begin 
      x02bai <= 32'b00111111100100111011111111001011;
      x02jyou <= 32'b00111110101010101000101110100110;
    end else if (wbdata[22:12] == 1501) begin 
      x02bai <= 32'b00111111100100111011010100100011;
      x02jyou <= 32'b00111110101010100111001100001101;
    end else if (wbdata[22:12] == 1502) begin 
      x02bai <= 32'b00111111100100111010101001111101;
      x02jyou <= 32'b00111110101010100101101001111010;
    end else if (wbdata[22:12] == 1503) begin 
      x02bai <= 32'b00111111100100111001111111011000;
      x02jyou <= 32'b00111110101010100100000111101100;
    end else if (wbdata[22:12] == 1504) begin 
      x02bai <= 32'b00111111100100111001010100110100;
      x02jyou <= 32'b00111110101010100010100101100001;
    end else if (wbdata[22:12] == 1505) begin 
      x02bai <= 32'b00111111100100111000101010010011;
      x02jyou <= 32'b00111110101010100001000011100000;
    end else if (wbdata[22:12] == 1506) begin 
      x02bai <= 32'b00111111100100110111111111110010;
      x02jyou <= 32'b00111110101010011111100001100000;
    end else if (wbdata[22:12] == 1507) begin 
      x02bai <= 32'b00111111100100110111010101010100;
      x02jyou <= 32'b00111110101010011101111111101000;
    end else if (wbdata[22:12] == 1508) begin 
      x02bai <= 32'b00111111100100110110101010110110;
      x02jyou <= 32'b00111110101010011100011101110011;
    end else if (wbdata[22:12] == 1509) begin 
      x02bai <= 32'b00111111100100110110000000011011;
      x02jyou <= 32'b00111110101010011010111100000110;
    end else if (wbdata[22:12] == 1510) begin 
      x02bai <= 32'b00111111100100110101010110000000;
      x02jyou <= 32'b00111110101010011001011010011011;
    end else if (wbdata[22:12] == 1511) begin 
      x02bai <= 32'b00111111100100110100101011101000;
      x02jyou <= 32'b00111110101010010111111000111001;
    end else if (wbdata[22:12] == 1512) begin 
      x02bai <= 32'b00111111100100110100000001010001;
      x02jyou <= 32'b00111110101010010110010111011010;
    end else if (wbdata[22:12] == 1513) begin 
      x02bai <= 32'b00111111100100110011010110111011;
      x02jyou <= 32'b00111110101010010100110110000000;
    end else if (wbdata[22:12] == 1514) begin 
      x02bai <= 32'b00111111100100110010101100100111;
      x02jyou <= 32'b00111110101010010011010100101100;
    end else if (wbdata[22:12] == 1515) begin 
      x02bai <= 32'b00111111100100110010000010010100;
      x02jyou <= 32'b00111110101010010001110011011100;
    end else if (wbdata[22:12] == 1516) begin 
      x02bai <= 32'b00111111100100110001011000000011;
      x02jyou <= 32'b00111110101010010000010010010011;
    end else if (wbdata[22:12] == 1517) begin 
      x02bai <= 32'b00111111100100110000101101110100;
      x02jyou <= 32'b00111110101010001110110001001111;
    end else if (wbdata[22:12] == 1518) begin 
      x02bai <= 32'b00111111100100110000000011100110;
      x02jyou <= 32'b00111110101010001101010000010000;
    end else if (wbdata[22:12] == 1519) begin 
      x02bai <= 32'b00111111100100101111011001011001;
      x02jyou <= 32'b00111110101010001011101111010101;
    end else if (wbdata[22:12] == 1520) begin 
      x02bai <= 32'b00111111100100101110101111001110;
      x02jyou <= 32'b00111110101010001010001110100000;
    end else if (wbdata[22:12] == 1521) begin 
      x02bai <= 32'b00111111100100101110000101000101;
      x02jyou <= 32'b00111110101010001000101101110010;
    end else if (wbdata[22:12] == 1522) begin 
      x02bai <= 32'b00111111100100101101011010111101;
      x02jyou <= 32'b00111110101010000111001101000111;
    end else if (wbdata[22:12] == 1523) begin 
      x02bai <= 32'b00111111100100101100110000110111;
      x02jyou <= 32'b00111110101010000101101100100011;
    end else if (wbdata[22:12] == 1524) begin 
      x02bai <= 32'b00111111100100101100000110110010;
      x02jyou <= 32'b00111110101010000100001100000011;
    end else if (wbdata[22:12] == 1525) begin 
      x02bai <= 32'b00111111100100101011011100101110;
      x02jyou <= 32'b00111110101010000010101011100111;
    end else if (wbdata[22:12] == 1526) begin 
      x02bai <= 32'b00111111100100101010110010101100;
      x02jyou <= 32'b00111110101010000001001011010001;
    end else if (wbdata[22:12] == 1527) begin 
      x02bai <= 32'b00111111100100101010001000101100;
      x02jyou <= 32'b00111110101001111111101011000010;
    end else if (wbdata[22:12] == 1528) begin 
      x02bai <= 32'b00111111100100101001011110101101;
      x02jyou <= 32'b00111110101001111110001010110110;
    end else if (wbdata[22:12] == 1529) begin 
      x02bai <= 32'b00111111100100101000110100101111;
      x02jyou <= 32'b00111110101001111100101010101111;
    end else if (wbdata[22:12] == 1530) begin 
      x02bai <= 32'b00111111100100101000001010110100;
      x02jyou <= 32'b00111110101001111011001010110000;
    end else if (wbdata[22:12] == 1531) begin 
      x02bai <= 32'b00111111100100100111100000111001;
      x02jyou <= 32'b00111110101001111001101010110011;
    end else if (wbdata[22:12] == 1532) begin 
      x02bai <= 32'b00111111100100100110110111000000;
      x02jyou <= 32'b00111110101001111000001010111100;
    end else if (wbdata[22:12] == 1533) begin 
      x02bai <= 32'b00111111100100100110001101001001;
      x02jyou <= 32'b00111110101001110110101011001100;
    end else if (wbdata[22:12] == 1534) begin 
      x02bai <= 32'b00111111100100100101100011010011;
      x02jyou <= 32'b00111110101001110101001011011111;
    end else if (wbdata[22:12] == 1535) begin 
      x02bai <= 32'b00111111100100100100111001011110;
      x02jyou <= 32'b00111110101001110011101011110110;
    end else if (wbdata[22:12] == 1536) begin 
      x02bai <= 32'b00111111100100100100001111101011;
      x02jyou <= 32'b00111110101001110010001100010100;
    end else if (wbdata[22:12] == 1537) begin 
      x02bai <= 32'b00111111100100100011100101111010;
      x02jyou <= 32'b00111110101001110000101100111000;
    end else if (wbdata[22:12] == 1538) begin 
      x02bai <= 32'b00111111100100100010111100001010;
      x02jyou <= 32'b00111110101001101111001101100000;
    end else if (wbdata[22:12] == 1539) begin 
      x02bai <= 32'b00111111100100100010010010011100;
      x02jyou <= 32'b00111110101001101101101110001110;
    end else if (wbdata[22:12] == 1540) begin 
      x02bai <= 32'b00111111100100100001101000101111;
      x02jyou <= 32'b00111110101001101100001111000001;
    end else if (wbdata[22:12] == 1541) begin 
      x02bai <= 32'b00111111100100100000111111000011;
      x02jyou <= 32'b00111110101001101010101111110111;
    end else if (wbdata[22:12] == 1542) begin 
      x02bai <= 32'b00111111100100100000010101011001;
      x02jyou <= 32'b00111110101001101001010000110011;
    end else if (wbdata[22:12] == 1543) begin 
      x02bai <= 32'b00111111100100011111101011110001;
      x02jyou <= 32'b00111110101001100111110001110110;
    end else if (wbdata[22:12] == 1544) begin 
      x02bai <= 32'b00111111100100011111000010001010;
      x02jyou <= 32'b00111110101001100110010010111101;
    end else if (wbdata[22:12] == 1545) begin 
      x02bai <= 32'b00111111100100011110011000100100;
      x02jyou <= 32'b00111110101001100100110100000111;
    end else if (wbdata[22:12] == 1546) begin 
      x02bai <= 32'b00111111100100011101101111000000;
      x02jyou <= 32'b00111110101001100011010101011000;
    end else if (wbdata[22:12] == 1547) begin 
      x02bai <= 32'b00111111100100011101000101011101;
      x02jyou <= 32'b00111110101001100001110110101101;
    end else if (wbdata[22:12] == 1548) begin 
      x02bai <= 32'b00111111100100011100011011111100;
      x02jyou <= 32'b00111110101001100000011000001000;
    end else if (wbdata[22:12] == 1549) begin 
      x02bai <= 32'b00111111100100011011110010011101;
      x02jyou <= 32'b00111110101001011110111001101010;
    end else if (wbdata[22:12] == 1550) begin 
      x02bai <= 32'b00111111100100011011001000111110;
      x02jyou <= 32'b00111110101001011101011011001101;
    end else if (wbdata[22:12] == 1551) begin 
      x02bai <= 32'b00111111100100011010011111100010;
      x02jyou <= 32'b00111110101001011011111100111000;
    end else if (wbdata[22:12] == 1552) begin 
      x02bai <= 32'b00111111100100011001110110000111;
      x02jyou <= 32'b00111110101001011010011110101000;
    end else if (wbdata[22:12] == 1553) begin 
      x02bai <= 32'b00111111100100011001001100101101;
      x02jyou <= 32'b00111110101001011001000000011011;
    end else if (wbdata[22:12] == 1554) begin 
      x02bai <= 32'b00111111100100011000100011010101;
      x02jyou <= 32'b00111110101001010111100010010101;
    end else if (wbdata[22:12] == 1555) begin 
      x02bai <= 32'b00111111100100010111111001111110;
      x02jyou <= 32'b00111110101001010110000100010010;
    end else if (wbdata[22:12] == 1556) begin 
      x02bai <= 32'b00111111100100010111010000101000;
      x02jyou <= 32'b00111110101001010100100110010100;
    end else if (wbdata[22:12] == 1557) begin 
      x02bai <= 32'b00111111100100010110100111010101;
      x02jyou <= 32'b00111110101001010011001000011110;
    end else if (wbdata[22:12] == 1558) begin 
      x02bai <= 32'b00111111100100010101111110000010;
      x02jyou <= 32'b00111110101001010001101010101010;
    end else if (wbdata[22:12] == 1559) begin 
      x02bai <= 32'b00111111100100010101010100110001;
      x02jyou <= 32'b00111110101001010000001100111100;
    end else if (wbdata[22:12] == 1560) begin 
      x02bai <= 32'b00111111100100010100101011100010;
      x02jyou <= 32'b00111110101001001110101111010100;
    end else if (wbdata[22:12] == 1561) begin 
      x02bai <= 32'b00111111100100010100000010010100;
      x02jyou <= 32'b00111110101001001101010001110000;
    end else if (wbdata[22:12] == 1562) begin 
      x02bai <= 32'b00111111100100010011011001000111;
      x02jyou <= 32'b00111110101001001011110100010000;
    end else if (wbdata[22:12] == 1563) begin 
      x02bai <= 32'b00111111100100010010101111111100;
      x02jyou <= 32'b00111110101001001010010110110110;
    end else if (wbdata[22:12] == 1564) begin 
      x02bai <= 32'b00111111100100010010000110110010;
      x02jyou <= 32'b00111110101001001000111001100000;
    end else if (wbdata[22:12] == 1565) begin 
      x02bai <= 32'b00111111100100010001011101101010;
      x02jyou <= 32'b00111110101001000111011100010000;
    end else if (wbdata[22:12] == 1566) begin 
      x02bai <= 32'b00111111100100010000110100100100;
      x02jyou <= 32'b00111110101001000101111111000111;
    end else if (wbdata[22:12] == 1567) begin 
      x02bai <= 32'b00111111100100010000001011011110;
      x02jyou <= 32'b00111110101001000100100001111111;
    end else if (wbdata[22:12] == 1568) begin 
      x02bai <= 32'b00111111100100001111100010011010;
      x02jyou <= 32'b00111110101001000011000100111101;
    end else if (wbdata[22:12] == 1569) begin 
      x02bai <= 32'b00111111100100001110111001011000;
      x02jyou <= 32'b00111110101001000001101000000010;
    end else if (wbdata[22:12] == 1570) begin 
      x02bai <= 32'b00111111100100001110010000010111;
      x02jyou <= 32'b00111110101001000000001011001010;
    end else if (wbdata[22:12] == 1571) begin 
      x02bai <= 32'b00111111100100001101100111011000;
      x02jyou <= 32'b00111110101000111110101110011001;
    end else if (wbdata[22:12] == 1572) begin 
      x02bai <= 32'b00111111100100001100111110011010;
      x02jyou <= 32'b00111110101000111101010001101011;
    end else if (wbdata[22:12] == 1573) begin 
      x02bai <= 32'b00111111100100001100010101011101;
      x02jyou <= 32'b00111110101000111011110101000010;
    end else if (wbdata[22:12] == 1574) begin 
      x02bai <= 32'b00111111100100001011101100100010;
      x02jyou <= 32'b00111110101000111010011000011110;
    end else if (wbdata[22:12] == 1575) begin 
      x02bai <= 32'b00111111100100001011000011101000;
      x02jyou <= 32'b00111110101000111000111011111110;
    end else if (wbdata[22:12] == 1576) begin 
      x02bai <= 32'b00111111100100001010011010110000;
      x02jyou <= 32'b00111110101000110111011111100101;
    end else if (wbdata[22:12] == 1577) begin 
      x02bai <= 32'b00111111100100001001110001111001;
      x02jyou <= 32'b00111110101000110110000011010000;
    end else if (wbdata[22:12] == 1578) begin 
      x02bai <= 32'b00111111100100001001001001000100;
      x02jyou <= 32'b00111110101000110100100111000000;
    end else if (wbdata[22:12] == 1579) begin 
      x02bai <= 32'b00111111100100001000100000010000;
      x02jyou <= 32'b00111110101000110011001010110101;
    end else if (wbdata[22:12] == 1580) begin 
      x02bai <= 32'b00111111100100000111110111011110;
      x02jyou <= 32'b00111110101000110001101110101111;
    end else if (wbdata[22:12] == 1581) begin 
      x02bai <= 32'b00111111100100000111001110101101;
      x02jyou <= 32'b00111110101000110000010010101110;
    end else if (wbdata[22:12] == 1582) begin 
      x02bai <= 32'b00111111100100000110100101111101;
      x02jyou <= 32'b00111110101000101110110110110000;
    end else if (wbdata[22:12] == 1583) begin 
      x02bai <= 32'b00111111100100000101111101001111;
      x02jyou <= 32'b00111110101000101101011010111001;
    end else if (wbdata[22:12] == 1584) begin 
      x02bai <= 32'b00111111100100000101010100100010;
      x02jyou <= 32'b00111110101000101011111111000101;
    end else if (wbdata[22:12] == 1585) begin 
      x02bai <= 32'b00111111100100000100101011110111;
      x02jyou <= 32'b00111110101000101010100011011000;
    end else if (wbdata[22:12] == 1586) begin 
      x02bai <= 32'b00111111100100000100000011001101;
      x02jyou <= 32'b00111110101000101001000111101110;
    end else if (wbdata[22:12] == 1587) begin 
      x02bai <= 32'b00111111100100000011011010100101;
      x02jyou <= 32'b00111110101000100111101100001011;
    end else if (wbdata[22:12] == 1588) begin 
      x02bai <= 32'b00111111100100000010110001111110;
      x02jyou <= 32'b00111110101000100110010000101011;
    end else if (wbdata[22:12] == 1589) begin 
      x02bai <= 32'b00111111100100000010001001011000;
      x02jyou <= 32'b00111110101000100100110101001111;
    end else if (wbdata[22:12] == 1590) begin 
      x02bai <= 32'b00111111100100000001100000110100;
      x02jyou <= 32'b00111110101000100011011001111010;
    end else if (wbdata[22:12] == 1591) begin 
      x02bai <= 32'b00111111100100000000111000010010;
      x02jyou <= 32'b00111110101000100001111110101010;
    end else if (wbdata[22:12] == 1592) begin 
      x02bai <= 32'b00111111100100000000001111110000;
      x02jyou <= 32'b00111110101000100000100011011100;
    end else if (wbdata[22:12] == 1593) begin 
      x02bai <= 32'b00111111100011111111100111010000;
      x02jyou <= 32'b00111110101000011111001000010100;
    end else if (wbdata[22:12] == 1594) begin 
      x02bai <= 32'b00111111100011111110111110110010;
      x02jyou <= 32'b00111110101000011101101101010011;
    end else if (wbdata[22:12] == 1595) begin 
      x02bai <= 32'b00111111100011111110010110010101;
      x02jyou <= 32'b00111110101000011100010010010101;
    end else if (wbdata[22:12] == 1596) begin 
      x02bai <= 32'b00111111100011111101101101111001;
      x02jyou <= 32'b00111110101000011010110111011011;
    end else if (wbdata[22:12] == 1597) begin 
      x02bai <= 32'b00111111100011111101000101011111;
      x02jyou <= 32'b00111110101000011001011100100111;
    end else if (wbdata[22:12] == 1598) begin 
      x02bai <= 32'b00111111100011111100011101000111;
      x02jyou <= 32'b00111110101000011000000001111001;
    end else if (wbdata[22:12] == 1599) begin 
      x02bai <= 32'b00111111100011111011110100101111;
      x02jyou <= 32'b00111110101000010110100111001101;
    end else if (wbdata[22:12] == 1600) begin 
      x02bai <= 32'b00111111100011111011001100011001;
      x02jyou <= 32'b00111110101000010101001100100110;
    end else if (wbdata[22:12] == 1601) begin 
      x02bai <= 32'b00111111100011111010100100000101;
      x02jyou <= 32'b00111110101000010011110010000110;
    end else if (wbdata[22:12] == 1602) begin 
      x02bai <= 32'b00111111100011111001111011110010;
      x02jyou <= 32'b00111110101000010010010111101010;
    end else if (wbdata[22:12] == 1603) begin 
      x02bai <= 32'b00111111100011111001010011100000;
      x02jyou <= 32'b00111110101000010000111101010010;
    end else if (wbdata[22:12] == 1604) begin 
      x02bai <= 32'b00111111100011111000101011010000;
      x02jyou <= 32'b00111110101000001111100010111111;
    end else if (wbdata[22:12] == 1605) begin 
      x02bai <= 32'b00111111100011111000000011000001;
      x02jyou <= 32'b00111110101000001110001000110001;
    end else if (wbdata[22:12] == 1606) begin 
      x02bai <= 32'b00111111100011110111011010110100;
      x02jyou <= 32'b00111110101000001100101110101000;
    end else if (wbdata[22:12] == 1607) begin 
      x02bai <= 32'b00111111100011110110110010101000;
      x02jyou <= 32'b00111110101000001011010100100100;
    end else if (wbdata[22:12] == 1608) begin 
      x02bai <= 32'b00111111100011110110001010011101;
      x02jyou <= 32'b00111110101000001001111010100011;
    end else if (wbdata[22:12] == 1609) begin 
      x02bai <= 32'b00111111100011110101100010010100;
      x02jyou <= 32'b00111110101000001000100000101000;
    end else if (wbdata[22:12] == 1610) begin 
      x02bai <= 32'b00111111100011110100111010001100;
      x02jyou <= 32'b00111110101000000111000110110001;
    end else if (wbdata[22:12] == 1611) begin 
      x02bai <= 32'b00111111100011110100010010000110;
      x02jyou <= 32'b00111110101000000101101101000000;
    end else if (wbdata[22:12] == 1612) begin 
      x02bai <= 32'b00111111100011110011101010000001;
      x02jyou <= 32'b00111110101000000100010011010011;
    end else if (wbdata[22:12] == 1613) begin 
      x02bai <= 32'b00111111100011110011000001111101;
      x02jyou <= 32'b00111110101000000010111001101010;
    end else if (wbdata[22:12] == 1614) begin 
      x02bai <= 32'b00111111100011110010011001111011;
      x02jyou <= 32'b00111110101000000001100000000110;
    end else if (wbdata[22:12] == 1615) begin 
      x02bai <= 32'b00111111100011110001110001111010;
      x02jyou <= 32'b00111110101000000000000110100111;
    end else if (wbdata[22:12] == 1616) begin 
      x02bai <= 32'b00111111100011110001001001111010;
      x02jyou <= 32'b00111110100111111110101101001011;
    end else if (wbdata[22:12] == 1617) begin 
      x02bai <= 32'b00111111100011110000100001111100;
      x02jyou <= 32'b00111110100111111101010011110110;
    end else if (wbdata[22:12] == 1618) begin 
      x02bai <= 32'b00111111100011101111111010000000;
      x02jyou <= 32'b00111110100111111011111010100110;
    end else if (wbdata[22:12] == 1619) begin 
      x02bai <= 32'b00111111100011101111010010000101;
      x02jyou <= 32'b00111110100111111010100001011010;
    end else if (wbdata[22:12] == 1620) begin 
      x02bai <= 32'b00111111100011101110101010001011;
      x02jyou <= 32'b00111110100111111001001000010010;
    end else if (wbdata[22:12] == 1621) begin 
      x02bai <= 32'b00111111100011101110000010010010;
      x02jyou <= 32'b00111110100111110111101111001110;
    end else if (wbdata[22:12] == 1622) begin 
      x02bai <= 32'b00111111100011101101011010011011;
      x02jyou <= 32'b00111110100111110110010110010000;
    end else if (wbdata[22:12] == 1623) begin 
      x02bai <= 32'b00111111100011101100110010100110;
      x02jyou <= 32'b00111110100111110100111101011000;
    end else if (wbdata[22:12] == 1624) begin 
      x02bai <= 32'b00111111100011101100001010110001;
      x02jyou <= 32'b00111110100111110011100100100001;
    end else if (wbdata[22:12] == 1625) begin 
      x02bai <= 32'b00111111100011101011100010111111;
      x02jyou <= 32'b00111110100111110010001011110010;
    end else if (wbdata[22:12] == 1626) begin 
      x02bai <= 32'b00111111100011101010111011001101;
      x02jyou <= 32'b00111110100111110000110011000110;
    end else if (wbdata[22:12] == 1627) begin 
      x02bai <= 32'b00111111100011101010010011011101;
      x02jyou <= 32'b00111110100111101111011010011111;
    end else if (wbdata[22:12] == 1628) begin 
      x02bai <= 32'b00111111100011101001101011101110;
      x02jyou <= 32'b00111110100111101110000001111100;
    end else if (wbdata[22:12] == 1629) begin 
      x02bai <= 32'b00111111100011101001000100000001;
      x02jyou <= 32'b00111110100111101100101001011110;
    end else if (wbdata[22:12] == 1630) begin 
      x02bai <= 32'b00111111100011101000011100010101;
      x02jyou <= 32'b00111110100111101011010001000101;
    end else if (wbdata[22:12] == 1631) begin 
      x02bai <= 32'b00111111100011100111110100101010;
      x02jyou <= 32'b00111110100111101001111000110000;
    end else if (wbdata[22:12] == 1632) begin 
      x02bai <= 32'b00111111100011100111001101000001;
      x02jyou <= 32'b00111110100111101000100000100000;
    end else if (wbdata[22:12] == 1633) begin 
      x02bai <= 32'b00111111100011100110100101011001;
      x02jyou <= 32'b00111110100111100111001000010100;
    end else if (wbdata[22:12] == 1634) begin 
      x02bai <= 32'b00111111100011100101111101110011;
      x02jyou <= 32'b00111110100111100101110000001110;
    end else if (wbdata[22:12] == 1635) begin 
      x02bai <= 32'b00111111100011100101010110001110;
      x02jyou <= 32'b00111110100111100100011000001100;
    end else if (wbdata[22:12] == 1636) begin 
      x02bai <= 32'b00111111100011100100101110101010;
      x02jyou <= 32'b00111110100111100011000000001110;
    end else if (wbdata[22:12] == 1637) begin 
      x02bai <= 32'b00111111100011100100000111001000;
      x02jyou <= 32'b00111110100111100001101000010110;
    end else if (wbdata[22:12] == 1638) begin 
      x02bai <= 32'b00111111100011100011011111100111;
      x02jyou <= 32'b00111110100111100000010000100001;
    end else if (wbdata[22:12] == 1639) begin 
      x02bai <= 32'b00111111100011100010111000000111;
      x02jyou <= 32'b00111110100111011110111000110000;
    end else if (wbdata[22:12] == 1640) begin 
      x02bai <= 32'b00111111100011100010010000101001;
      x02jyou <= 32'b00111110100111011101100001000101;
    end else if (wbdata[22:12] == 1641) begin 
      x02bai <= 32'b00111111100011100001101001001100;
      x02jyou <= 32'b00111110100111011100001001011110;
    end else if (wbdata[22:12] == 1642) begin 
      x02bai <= 32'b00111111100011100001000001110001;
      x02jyou <= 32'b00111110100111011010110001111101;
    end else if (wbdata[22:12] == 1643) begin 
      x02bai <= 32'b00111111100011100000011010010111;
      x02jyou <= 32'b00111110100111011001011010011111;
    end else if (wbdata[22:12] == 1644) begin 
      x02bai <= 32'b00111111100011011111110010111110;
      x02jyou <= 32'b00111110100111011000000011000110;
    end else if (wbdata[22:12] == 1645) begin 
      x02bai <= 32'b00111111100011011111001011100111;
      x02jyou <= 32'b00111110100111010110101011110010;
    end else if (wbdata[22:12] == 1646) begin 
      x02bai <= 32'b00111111100011011110100100010001;
      x02jyou <= 32'b00111110100111010101010100100010;
    end else if (wbdata[22:12] == 1647) begin 
      x02bai <= 32'b00111111100011011101111100111100;
      x02jyou <= 32'b00111110100111010011111101010110;
    end else if (wbdata[22:12] == 1648) begin 
      x02bai <= 32'b00111111100011011101010101101001;
      x02jyou <= 32'b00111110100111010010100110001111;
    end else if (wbdata[22:12] == 1649) begin 
      x02bai <= 32'b00111111100011011100101110010111;
      x02jyou <= 32'b00111110100111010001001111001100;
    end else if (wbdata[22:12] == 1650) begin 
      x02bai <= 32'b00111111100011011100000111000110;
      x02jyou <= 32'b00111110100111001111111000001110;
    end else if (wbdata[22:12] == 1651) begin 
      x02bai <= 32'b00111111100011011011011111110111;
      x02jyou <= 32'b00111110100111001110100001010101;
    end else if (wbdata[22:12] == 1652) begin 
      x02bai <= 32'b00111111100011011010111000101001;
      x02jyou <= 32'b00111110100111001101001010011111;
    end else if (wbdata[22:12] == 1653) begin 
      x02bai <= 32'b00111111100011011010010001011101;
      x02jyou <= 32'b00111110100111001011110011110000;
    end else if (wbdata[22:12] == 1654) begin 
      x02bai <= 32'b00111111100011011001101010010010;
      x02jyou <= 32'b00111110100111001010011101000100;
    end else if (wbdata[22:12] == 1655) begin 
      x02bai <= 32'b00111111100011011001000011001000;
      x02jyou <= 32'b00111110100111001001000110011100;
    end else if (wbdata[22:12] == 1656) begin 
      x02bai <= 32'b00111111100011011000011011111111;
      x02jyou <= 32'b00111110100111000111101111111000;
    end else if (wbdata[22:12] == 1657) begin 
      x02bai <= 32'b00111111100011010111110100111000;
      x02jyou <= 32'b00111110100111000110011001011010;
    end else if (wbdata[22:12] == 1658) begin 
      x02bai <= 32'b00111111100011010111001101110011;
      x02jyou <= 32'b00111110100111000101000011000001;
    end else if (wbdata[22:12] == 1659) begin 
      x02bai <= 32'b00111111100011010110100110101110;
      x02jyou <= 32'b00111110100111000011101100101011;
    end else if (wbdata[22:12] == 1660) begin 
      x02bai <= 32'b00111111100011010101111111101011;
      x02jyou <= 32'b00111110100111000010010110011010;
    end else if (wbdata[22:12] == 1661) begin 
      x02bai <= 32'b00111111100011010101011000101010;
      x02jyou <= 32'b00111110100111000001000000001111;
    end else if (wbdata[22:12] == 1662) begin 
      x02bai <= 32'b00111111100011010100110001101001;
      x02jyou <= 32'b00111110100110111111101010000101;
    end else if (wbdata[22:12] == 1663) begin 
      x02bai <= 32'b00111111100011010100001010101010;
      x02jyou <= 32'b00111110100110111110010100000001;
    end else if (wbdata[22:12] == 1664) begin 
      x02bai <= 32'b00111111100011010011100011101101;
      x02jyou <= 32'b00111110100110111100111110000011;
    end else if (wbdata[22:12] == 1665) begin 
      x02bai <= 32'b00111111100011010010111100110000;
      x02jyou <= 32'b00111110100110111011101000000111;
    end else if (wbdata[22:12] == 1666) begin 
      x02bai <= 32'b00111111100011010010010101110101;
      x02jyou <= 32'b00111110100110111010010010010001;
    end else if (wbdata[22:12] == 1667) begin 
      x02bai <= 32'b00111111100011010001101110111100;
      x02jyou <= 32'b00111110100110111000111100100000;
    end else if (wbdata[22:12] == 1668) begin 
      x02bai <= 32'b00111111100011010001001000000011;
      x02jyou <= 32'b00111110100110110111100110110001;
    end else if (wbdata[22:12] == 1669) begin 
      x02bai <= 32'b00111111100011010000100001001100;
      x02jyou <= 32'b00111110100110110110010001001000;
    end else if (wbdata[22:12] == 1670) begin 
      x02bai <= 32'b00111111100011001111111010010111;
      x02jyou <= 32'b00111110100110110100111011100101;
    end else if (wbdata[22:12] == 1671) begin 
      x02bai <= 32'b00111111100011001111010011100011;
      x02jyou <= 32'b00111110100110110011100110000101;
    end else if (wbdata[22:12] == 1672) begin 
      x02bai <= 32'b00111111100011001110101100110000;
      x02jyou <= 32'b00111110100110110010010000101001;
    end else if (wbdata[22:12] == 1673) begin 
      x02bai <= 32'b00111111100011001110000101111110;
      x02jyou <= 32'b00111110100110110000111011010001;
    end else if (wbdata[22:12] == 1674) begin 
      x02bai <= 32'b00111111100011001101011111001110;
      x02jyou <= 32'b00111110100110101111100101111110;
    end else if (wbdata[22:12] == 1675) begin 
      x02bai <= 32'b00111111100011001100111000011111;
      x02jyou <= 32'b00111110100110101110010000110000;
    end else if (wbdata[22:12] == 1676) begin 
      x02bai <= 32'b00111111100011001100010001110001;
      x02jyou <= 32'b00111110100110101100111011100101;
    end else if (wbdata[22:12] == 1677) begin 
      x02bai <= 32'b00111111100011001011101011000101;
      x02jyou <= 32'b00111110100110101011100110011111;
    end else if (wbdata[22:12] == 1678) begin 
      x02bai <= 32'b00111111100011001011000100011010;
      x02jyou <= 32'b00111110100110101010010001011110;
    end else if (wbdata[22:12] == 1679) begin 
      x02bai <= 32'b00111111100011001010011101110000;
      x02jyou <= 32'b00111110100110101000111100100000;
    end else if (wbdata[22:12] == 1680) begin 
      x02bai <= 32'b00111111100011001001110111001000;
      x02jyou <= 32'b00111110100110100111100111101000;
    end else if (wbdata[22:12] == 1681) begin 
      x02bai <= 32'b00111111100011001001010000100001;
      x02jyou <= 32'b00111110100110100110010010110100;
    end else if (wbdata[22:12] == 1682) begin 
      x02bai <= 32'b00111111100011001000101001111100;
      x02jyou <= 32'b00111110100110100100111110000101;
    end else if (wbdata[22:12] == 1683) begin 
      x02bai <= 32'b00111111100011001000000011010111;
      x02jyou <= 32'b00111110100110100011101001011000;
    end else if (wbdata[22:12] == 1684) begin 
      x02bai <= 32'b00111111100011000111011100110100;
      x02jyou <= 32'b00111110100110100010010100110001;
    end else if (wbdata[22:12] == 1685) begin 
      x02bai <= 32'b00111111100011000110110110010011;
      x02jyou <= 32'b00111110100110100001000000001111;
    end else if (wbdata[22:12] == 1686) begin 
      x02bai <= 32'b00111111100011000110001111110010;
      x02jyou <= 32'b00111110100110011111101011101111;
    end else if (wbdata[22:12] == 1687) begin 
      x02bai <= 32'b00111111100011000101101001010011;
      x02jyou <= 32'b00111110100110011110010111010101;
    end else if (wbdata[22:12] == 1688) begin 
      x02bai <= 32'b00111111100011000101000010110110;
      x02jyou <= 32'b00111110100110011101000011000001;
    end else if (wbdata[22:12] == 1689) begin 
      x02bai <= 32'b00111111100011000100011100011001;
      x02jyou <= 32'b00111110100110011011101110101110;
    end else if (wbdata[22:12] == 1690) begin 
      x02bai <= 32'b00111111100011000011110101111110;
      x02jyou <= 32'b00111110100110011010011010100001;
    end else if (wbdata[22:12] == 1691) begin 
      x02bai <= 32'b00111111100011000011001111100100;
      x02jyou <= 32'b00111110100110011001000110011000;
    end else if (wbdata[22:12] == 1692) begin 
      x02bai <= 32'b00111111100011000010101001001100;
      x02jyou <= 32'b00111110100110010111110010010100;
    end else if (wbdata[22:12] == 1693) begin 
      x02bai <= 32'b00111111100011000010000010110101;
      x02jyou <= 32'b00111110100110010110011110010100;
    end else if (wbdata[22:12] == 1694) begin 
      x02bai <= 32'b00111111100011000001011100011111;
      x02jyou <= 32'b00111110100110010101001010011000;
    end else if (wbdata[22:12] == 1695) begin 
      x02bai <= 32'b00111111100011000000110110001010;
      x02jyou <= 32'b00111110100110010011110110011111;
    end else if (wbdata[22:12] == 1696) begin 
      x02bai <= 32'b00111111100011000000001111110111;
      x02jyou <= 32'b00111110100110010010100010101100;
    end else if (wbdata[22:12] == 1697) begin 
      x02bai <= 32'b00111111100010111111101001100101;
      x02jyou <= 32'b00111110100110010001001110111101;
    end else if (wbdata[22:12] == 1698) begin 
      x02bai <= 32'b00111111100010111111000011010101;
      x02jyou <= 32'b00111110100110001111111011010100;
    end else if (wbdata[22:12] == 1699) begin 
      x02bai <= 32'b00111111100010111110011101000110;
      x02jyou <= 32'b00111110100110001110100111101110;
    end else if (wbdata[22:12] == 1700) begin 
      x02bai <= 32'b00111111100010111101110110111000;
      x02jyou <= 32'b00111110100110001101010100001100;
    end else if (wbdata[22:12] == 1701) begin 
      x02bai <= 32'b00111111100010111101010000101011;
      x02jyou <= 32'b00111110100110001100000000101101;
    end else if (wbdata[22:12] == 1702) begin 
      x02bai <= 32'b00111111100010111100101010100000;
      x02jyou <= 32'b00111110100110001010101101010100;
    end else if (wbdata[22:12] == 1703) begin 
      x02bai <= 32'b00111111100010111100000100010101;
      x02jyou <= 32'b00111110100110001001011001111101;
    end else if (wbdata[22:12] == 1704) begin 
      x02bai <= 32'b00111111100010111011011110001101;
      x02jyou <= 32'b00111110100110001000000110101101;
    end else if (wbdata[22:12] == 1705) begin 
      x02bai <= 32'b00111111100010111010111000000101;
      x02jyou <= 32'b00111110100110000110110011011111;
    end else if (wbdata[22:12] == 1706) begin 
      x02bai <= 32'b00111111100010111010010001111111;
      x02jyou <= 32'b00111110100110000101100000010111;
    end else if (wbdata[22:12] == 1707) begin 
      x02bai <= 32'b00111111100010111001101011111010;
      x02jyou <= 32'b00111110100110000100001101010011;
    end else if (wbdata[22:12] == 1708) begin 
      x02bai <= 32'b00111111100010111001000101110111;
      x02jyou <= 32'b00111110100110000010111010010100;
    end else if (wbdata[22:12] == 1709) begin 
      x02bai <= 32'b00111111100010111000011111110100;
      x02jyou <= 32'b00111110100110000001100111010110;
    end else if (wbdata[22:12] == 1710) begin 
      x02bai <= 32'b00111111100010110111111001110011;
      x02jyou <= 32'b00111110100110000000010100011111;
    end else if (wbdata[22:12] == 1711) begin 
      x02bai <= 32'b00111111100010110111010011110100;
      x02jyou <= 32'b00111110100101111111000001101101;
    end else if (wbdata[22:12] == 1712) begin 
      x02bai <= 32'b00111111100010110110101101110101;
      x02jyou <= 32'b00111110100101111101101110111100;
    end else if (wbdata[22:12] == 1713) begin 
      x02bai <= 32'b00111111100010110110000111111000;
      x02jyou <= 32'b00111110100101111100011100010010;
    end else if (wbdata[22:12] == 1714) begin 
      x02bai <= 32'b00111111100010110101100001111101;
      x02jyou <= 32'b00111110100101111011001001101101;
    end else if (wbdata[22:12] == 1715) begin 
      x02bai <= 32'b00111111100010110100111100000010;
      x02jyou <= 32'b00111110100101111001110111001001;
    end else if (wbdata[22:12] == 1716) begin 
      x02bai <= 32'b00111111100010110100010110001001;
      x02jyou <= 32'b00111110100101111000100100101011;
    end else if (wbdata[22:12] == 1717) begin 
      x02bai <= 32'b00111111100010110011110000010001;
      x02jyou <= 32'b00111110100101110111010010010001;
    end else if (wbdata[22:12] == 1718) begin 
      x02bai <= 32'b00111111100010110011001010011010;
      x02jyou <= 32'b00111110100101110101111111111010;
    end else if (wbdata[22:12] == 1719) begin 
      x02bai <= 32'b00111111100010110010100100100101;
      x02jyou <= 32'b00111110100101110100101101101010;
    end else if (wbdata[22:12] == 1720) begin 
      x02bai <= 32'b00111111100010110001111110110001;
      x02jyou <= 32'b00111110100101110011011011011100;
    end else if (wbdata[22:12] == 1721) begin 
      x02bai <= 32'b00111111100010110001011000111110;
      x02jyou <= 32'b00111110100101110010001001010011;
    end else if (wbdata[22:12] == 1722) begin 
      x02bai <= 32'b00111111100010110000110011001101;
      x02jyou <= 32'b00111110100101110000110111001111;
    end else if (wbdata[22:12] == 1723) begin 
      x02bai <= 32'b00111111100010110000001101011100;
      x02jyou <= 32'b00111110100101101111100101001100;
    end else if (wbdata[22:12] == 1724) begin 
      x02bai <= 32'b00111111100010101111100111101101;
      x02jyou <= 32'b00111110100101101110010011001111;
    end else if (wbdata[22:12] == 1725) begin 
      x02bai <= 32'b00111111100010101111000010000000;
      x02jyou <= 32'b00111110100101101101000001011000;
    end else if (wbdata[22:12] == 1726) begin 
      x02bai <= 32'b00111111100010101110011100010011;
      x02jyou <= 32'b00111110100101101011101111100010;
    end else if (wbdata[22:12] == 1727) begin 
      x02bai <= 32'b00111111100010101101110110101000;
      x02jyou <= 32'b00111110100101101010011101110010;
    end else if (wbdata[22:12] == 1728) begin 
      x02bai <= 32'b00111111100010101101010000111110;
      x02jyou <= 32'b00111110100101101001001100000110;
    end else if (wbdata[22:12] == 1729) begin 
      x02bai <= 32'b00111111100010101100101011010110;
      x02jyou <= 32'b00111110100101100111111010011111;
    end else if (wbdata[22:12] == 1730) begin 
      x02bai <= 32'b00111111100010101100000101101111;
      x02jyou <= 32'b00111110100101100110101000111100;
    end else if (wbdata[22:12] == 1731) begin 
      x02bai <= 32'b00111111100010101011100000001001;
      x02jyou <= 32'b00111110100101100101010111011100;
    end else if (wbdata[22:12] == 1732) begin 
      x02bai <= 32'b00111111100010101010111010100100;
      x02jyou <= 32'b00111110100101100100000110000000;
    end else if (wbdata[22:12] == 1733) begin 
      x02bai <= 32'b00111111100010101010010101000000;
      x02jyou <= 32'b00111110100101100010110100100111;
    end else if (wbdata[22:12] == 1734) begin 
      x02bai <= 32'b00111111100010101001101111011110;
      x02jyou <= 32'b00111110100101100001100011010100;
    end else if (wbdata[22:12] == 1735) begin 
      x02bai <= 32'b00111111100010101001001001111101;
      x02jyou <= 32'b00111110100101100000010010000101;
    end else if (wbdata[22:12] == 1736) begin 
      x02bai <= 32'b00111111100010101000100100011110;
      x02jyou <= 32'b00111110100101011111000000111100;
    end else if (wbdata[22:12] == 1737) begin 
      x02bai <= 32'b00111111100010100111111110111111;
      x02jyou <= 32'b00111110100101011101101111110011;
    end else if (wbdata[22:12] == 1738) begin 
      x02bai <= 32'b00111111100010100111011001100010;
      x02jyou <= 32'b00111110100101011100011110110001;
    end else if (wbdata[22:12] == 1739) begin 
      x02bai <= 32'b00111111100010100110110100000110;
      x02jyou <= 32'b00111110100101011011001101110010;
    end else if (wbdata[22:12] == 1740) begin 
      x02bai <= 32'b00111111100010100110001110101100;
      x02jyou <= 32'b00111110100101011001111100111000;
    end else if (wbdata[22:12] == 1741) begin 
      x02bai <= 32'b00111111100010100101101001010010;
      x02jyou <= 32'b00111110100101011000101100000001;
    end else if (wbdata[22:12] == 1742) begin 
      x02bai <= 32'b00111111100010100101000011111010;
      x02jyou <= 32'b00111110100101010111011011001110;
    end else if (wbdata[22:12] == 1743) begin 
      x02bai <= 32'b00111111100010100100011110100100;
      x02jyou <= 32'b00111110100101010110001010100010;
    end else if (wbdata[22:12] == 1744) begin 
      x02bai <= 32'b00111111100010100011111001001110;
      x02jyou <= 32'b00111110100101010100111001110111;
    end else if (wbdata[22:12] == 1745) begin 
      x02bai <= 32'b00111111100010100011010011111010;
      x02jyou <= 32'b00111110100101010011101001010001;
    end else if (wbdata[22:12] == 1746) begin 
      x02bai <= 32'b00111111100010100010101110100111;
      x02jyou <= 32'b00111110100101010010011000101111;
    end else if (wbdata[22:12] == 1747) begin 
      x02bai <= 32'b00111111100010100010001001010101;
      x02jyou <= 32'b00111110100101010001001000010000;
    end else if (wbdata[22:12] == 1748) begin 
      x02bai <= 32'b00111111100010100001100100000100;
      x02jyou <= 32'b00111110100101001111110111110110;
    end else if (wbdata[22:12] == 1749) begin 
      x02bai <= 32'b00111111100010100000111110110101;
      x02jyou <= 32'b00111110100101001110100111100000;
    end else if (wbdata[22:12] == 1750) begin 
      x02bai <= 32'b00111111100010100000011001100111;
      x02jyou <= 32'b00111110100101001101010111001110;
    end else if (wbdata[22:12] == 1751) begin 
      x02bai <= 32'b00111111100010011111110100011010;
      x02jyou <= 32'b00111110100101001100000111000000;
    end else if (wbdata[22:12] == 1752) begin 
      x02bai <= 32'b00111111100010011111001111001111;
      x02jyou <= 32'b00111110100101001010110110111000;
    end else if (wbdata[22:12] == 1753) begin 
      x02bai <= 32'b00111111100010011110101010000101;
      x02jyou <= 32'b00111110100101001001100110110010;
    end else if (wbdata[22:12] == 1754) begin 
      x02bai <= 32'b00111111100010011110000100111100;
      x02jyou <= 32'b00111110100101001000010110110001;
    end else if (wbdata[22:12] == 1755) begin 
      x02bai <= 32'b00111111100010011101011111110100;
      x02jyou <= 32'b00111110100101000111000110110011;
    end else if (wbdata[22:12] == 1756) begin 
      x02bai <= 32'b00111111100010011100111010101110;
      x02jyou <= 32'b00111110100101000101110110111010;
    end else if (wbdata[22:12] == 1757) begin 
      x02bai <= 32'b00111111100010011100010101101000;
      x02jyou <= 32'b00111110100101000100100111000011;
    end else if (wbdata[22:12] == 1758) begin 
      x02bai <= 32'b00111111100010011011110000100100;
      x02jyou <= 32'b00111110100101000011010111010010;
    end else if (wbdata[22:12] == 1759) begin 
      x02bai <= 32'b00111111100010011011001011100010;
      x02jyou <= 32'b00111110100101000010000111100110;
    end else if (wbdata[22:12] == 1760) begin 
      x02bai <= 32'b00111111100010011010100110100000;
      x02jyou <= 32'b00111110100101000000110111111011;
    end else if (wbdata[22:12] == 1761) begin 
      x02bai <= 32'b00111111100010011010000001100000;
      x02jyou <= 32'b00111110100100111111101000010110;
    end else if (wbdata[22:12] == 1762) begin 
      x02bai <= 32'b00111111100010011001011100100001;
      x02jyou <= 32'b00111110100100111110011000110101;
    end else if (wbdata[22:12] == 1763) begin 
      x02bai <= 32'b00111111100010011000110111100011;
      x02jyou <= 32'b00111110100100111101001001010111;
    end else if (wbdata[22:12] == 1764) begin 
      x02bai <= 32'b00111111100010011000010010100111;
      x02jyou <= 32'b00111110100100111011111001111111;
    end else if (wbdata[22:12] == 1765) begin 
      x02bai <= 32'b00111111100010010111101101101011;
      x02jyou <= 32'b00111110100100111010101010101000;
    end else if (wbdata[22:12] == 1766) begin 
      x02bai <= 32'b00111111100010010111001000110001;
      x02jyou <= 32'b00111110100100111001011011010111;
    end else if (wbdata[22:12] == 1767) begin 
      x02bai <= 32'b00111111100010010110100011111000;
      x02jyou <= 32'b00111110100100111000001100001001;
    end else if (wbdata[22:12] == 1768) begin 
      x02bai <= 32'b00111111100010010101111111000001;
      x02jyou <= 32'b00111110100100110110111101000001;
    end else if (wbdata[22:12] == 1769) begin 
      x02bai <= 32'b00111111100010010101011010001010;
      x02jyou <= 32'b00111110100100110101101101111010;
    end else if (wbdata[22:12] == 1770) begin 
      x02bai <= 32'b00111111100010010100110101010101;
      x02jyou <= 32'b00111110100100110100011110111001;
    end else if (wbdata[22:12] == 1771) begin 
      x02bai <= 32'b00111111100010010100010000100010;
      x02jyou <= 32'b00111110100100110011001111111101;
    end else if (wbdata[22:12] == 1772) begin 
      x02bai <= 32'b00111111100010010011101011101111;
      x02jyou <= 32'b00111110100100110010000001000011;
    end else if (wbdata[22:12] == 1773) begin 
      x02bai <= 32'b00111111100010010011000110111101;
      x02jyou <= 32'b00111110100100110000110010001100;
    end else if (wbdata[22:12] == 1774) begin 
      x02bai <= 32'b00111111100010010010100010001101;
      x02jyou <= 32'b00111110100100101111100011011011;
    end else if (wbdata[22:12] == 1775) begin 
      x02bai <= 32'b00111111100010010001111101011110;
      x02jyou <= 32'b00111110100100101110010100101101;
    end else if (wbdata[22:12] == 1776) begin 
      x02bai <= 32'b00111111100010010001011000110001;
      x02jyou <= 32'b00111110100100101101000110000101;
    end else if (wbdata[22:12] == 1777) begin 
      x02bai <= 32'b00111111100010010000110100000100;
      x02jyou <= 32'b00111110100100101011110111011110;
    end else if (wbdata[22:12] == 1778) begin 
      x02bai <= 32'b00111111100010010000001111011001;
      x02jyou <= 32'b00111110100100101010101000111101;
    end else if (wbdata[22:12] == 1779) begin 
      x02bai <= 32'b00111111100010001111101010101111;
      x02jyou <= 32'b00111110100100101001011010011111;
    end else if (wbdata[22:12] == 1780) begin 
      x02bai <= 32'b00111111100010001111000110000110;
      x02jyou <= 32'b00111110100100101000001100000100;
    end else if (wbdata[22:12] == 1781) begin 
      x02bai <= 32'b00111111100010001110100001011111;
      x02jyou <= 32'b00111110100100100110111101110000;
    end else if (wbdata[22:12] == 1782) begin 
      x02bai <= 32'b00111111100010001101111100111000;
      x02jyou <= 32'b00111110100100100101101111011100;
    end else if (wbdata[22:12] == 1783) begin 
      x02bai <= 32'b00111111100010001101011000010011;
      x02jyou <= 32'b00111110100100100100100001001110;
    end else if (wbdata[22:12] == 1784) begin 
      x02bai <= 32'b00111111100010001100110011101111;
      x02jyou <= 32'b00111110100100100011010011000100;
    end else if (wbdata[22:12] == 1785) begin 
      x02bai <= 32'b00111111100010001100001111001100;
      x02jyou <= 32'b00111110100100100010000100111101;
    end else if (wbdata[22:12] == 1786) begin 
      x02bai <= 32'b00111111100010001011101010101011;
      x02jyou <= 32'b00111110100100100000110110111100;
    end else if (wbdata[22:12] == 1787) begin 
      x02bai <= 32'b00111111100010001011000110001011;
      x02jyou <= 32'b00111110100100011111101000111110;
    end else if (wbdata[22:12] == 1788) begin 
      x02bai <= 32'b00111111100010001010100001101100;
      x02jyou <= 32'b00111110100100011110011011000011;
    end else if (wbdata[22:12] == 1789) begin 
      x02bai <= 32'b00111111100010001001111101001110;
      x02jyou <= 32'b00111110100100011101001101001100;
    end else if (wbdata[22:12] == 1790) begin 
      x02bai <= 32'b00111111100010001001011000110001;
      x02jyou <= 32'b00111110100100011011111111011000;
    end else if (wbdata[22:12] == 1791) begin 
      x02bai <= 32'b00111111100010001000110100010110;
      x02jyou <= 32'b00111110100100011010110001101010;
    end else if (wbdata[22:12] == 1792) begin 
      x02bai <= 32'b00111111100010001000001111111100;
      x02jyou <= 32'b00111110100100011001100100000000;
    end else if (wbdata[22:12] == 1793) begin 
      x02bai <= 32'b00111111100010000111101011100011;
      x02jyou <= 32'b00111110100100011000010110011000;
    end else if (wbdata[22:12] == 1794) begin 
      x02bai <= 32'b00111111100010000111000111001011;
      x02jyou <= 32'b00111110100100010111001000110101;
    end else if (wbdata[22:12] == 1795) begin 
      x02bai <= 32'b00111111100010000110100010110101;
      x02jyou <= 32'b00111110100100010101111011010110;
    end else if (wbdata[22:12] == 1796) begin 
      x02bai <= 32'b00111111100010000101111110011111;
      x02jyou <= 32'b00111110100100010100101101111001;
    end else if (wbdata[22:12] == 1797) begin 
      x02bai <= 32'b00111111100010000101011010001011;
      x02jyou <= 32'b00111110100100010011100000100010;
    end else if (wbdata[22:12] == 1798) begin 
      x02bai <= 32'b00111111100010000100110101111000;
      x02jyou <= 32'b00111110100100010010010011001110;
    end else if (wbdata[22:12] == 1799) begin 
      x02bai <= 32'b00111111100010000100010001100110;
      x02jyou <= 32'b00111110100100010001000101111101;
    end else if (wbdata[22:12] == 1800) begin 
      x02bai <= 32'b00111111100010000011101101010110;
      x02jyou <= 32'b00111110100100001111111000110010;
    end else if (wbdata[22:12] == 1801) begin 
      x02bai <= 32'b00111111100010000011001001000111;
      x02jyou <= 32'b00111110100100001110101011101011;
    end else if (wbdata[22:12] == 1802) begin 
      x02bai <= 32'b00111111100010000010100100111001;
      x02jyou <= 32'b00111110100100001101011110100110;
    end else if (wbdata[22:12] == 1803) begin 
      x02bai <= 32'b00111111100010000010000000101100;
      x02jyou <= 32'b00111110100100001100010001100110;
    end else if (wbdata[22:12] == 1804) begin 
      x02bai <= 32'b00111111100010000001011100100000;
      x02jyou <= 32'b00111110100100001011000100101000;
    end else if (wbdata[22:12] == 1805) begin 
      x02bai <= 32'b00111111100010000000111000010110;
      x02jyou <= 32'b00111110100100001001110111110000;
    end else if (wbdata[22:12] == 1806) begin 
      x02bai <= 32'b00111111100010000000010100001100;
      x02jyou <= 32'b00111110100100001000101010111010;
    end else if (wbdata[22:12] == 1807) begin 
      x02bai <= 32'b00111111100001111111110000000100;
      x02jyou <= 32'b00111110100100000111011110001001;
    end else if (wbdata[22:12] == 1808) begin 
      x02bai <= 32'b00111111100001111111001011111101;
      x02jyou <= 32'b00111110100100000110010001011011;
    end else if (wbdata[22:12] == 1809) begin 
      x02bai <= 32'b00111111100001111110100111111000;
      x02jyou <= 32'b00111110100100000101000100110011;
    end else if (wbdata[22:12] == 1810) begin 
      x02bai <= 32'b00111111100001111110000011110011;
      x02jyou <= 32'b00111110100100000011111000001100;
    end else if (wbdata[22:12] == 1811) begin 
      x02bai <= 32'b00111111100001111101011111110000;
      x02jyou <= 32'b00111110100100000010101011101011;
    end else if (wbdata[22:12] == 1812) begin 
      x02bai <= 32'b00111111100001111100111011101110;
      x02jyou <= 32'b00111110100100000001011111001101;
    end else if (wbdata[22:12] == 1813) begin 
      x02bai <= 32'b00111111100001111100010111101101;
      x02jyou <= 32'b00111110100100000000010010110010;
    end else if (wbdata[22:12] == 1814) begin 
      x02bai <= 32'b00111111100001111011110011101101;
      x02jyou <= 32'b00111110100011111111000110011011;
    end else if (wbdata[22:12] == 1815) begin 
      x02bai <= 32'b00111111100001111011001111101111;
      x02jyou <= 32'b00111110100011111101111010001001;
    end else if (wbdata[22:12] == 1816) begin 
      x02bai <= 32'b00111111100001111010101011110001;
      x02jyou <= 32'b00111110100011111100101101111001;
    end else if (wbdata[22:12] == 1817) begin 
      x02bai <= 32'b00111111100001111010000111110101;
      x02jyou <= 32'b00111110100011111011100001101110;
    end else if (wbdata[22:12] == 1818) begin 
      x02bai <= 32'b00111111100001111001100011111010;
      x02jyou <= 32'b00111110100011111010010101100110;
    end else if (wbdata[22:12] == 1819) begin 
      x02bai <= 32'b00111111100001111001000000000001;
      x02jyou <= 32'b00111110100011111001001001100100;
    end else if (wbdata[22:12] == 1820) begin 
      x02bai <= 32'b00111111100001111000011100001000;
      x02jyou <= 32'b00111110100011110111111101100011;
    end else if (wbdata[22:12] == 1821) begin 
      x02bai <= 32'b00111111100001110111111000010001;
      x02jyou <= 32'b00111110100011110110110001101000;
    end else if (wbdata[22:12] == 1822) begin 
      x02bai <= 32'b00111111100001110111010100011011;
      x02jyou <= 32'b00111110100011110101100101110000;
    end else if (wbdata[22:12] == 1823) begin 
      x02bai <= 32'b00111111100001110110110000100110;
      x02jyou <= 32'b00111110100011110100011001111100;
    end else if (wbdata[22:12] == 1824) begin 
      x02bai <= 32'b00111111100001110110001100110010;
      x02jyou <= 32'b00111110100011110011001110001010;
    end else if (wbdata[22:12] == 1825) begin 
      x02bai <= 32'b00111111100001110101101000111111;
      x02jyou <= 32'b00111110100011110010000010011101;
    end else if (wbdata[22:12] == 1826) begin 
      x02bai <= 32'b00111111100001110101000101001110;
      x02jyou <= 32'b00111110100011110000110110110100;
    end else if (wbdata[22:12] == 1827) begin 
      x02bai <= 32'b00111111100001110100100001011101;
      x02jyou <= 32'b00111110100011101111101011001101;
    end else if (wbdata[22:12] == 1828) begin 
      x02bai <= 32'b00111111100001110011111101101110;
      x02jyou <= 32'b00111110100011101110011111101011;
    end else if (wbdata[22:12] == 1829) begin 
      x02bai <= 32'b00111111100001110011011010000000;
      x02jyou <= 32'b00111110100011101101010100001101;
    end else if (wbdata[22:12] == 1830) begin 
      x02bai <= 32'b00111111100001110010110110010100;
      x02jyou <= 32'b00111110100011101100001000110100;
    end else if (wbdata[22:12] == 1831) begin 
      x02bai <= 32'b00111111100001110010010010101000;
      x02jyou <= 32'b00111110100011101010111101011101;
    end else if (wbdata[22:12] == 1832) begin 
      x02bai <= 32'b00111111100001110001101110111110;
      x02jyou <= 32'b00111110100011101001110010001011;
    end else if (wbdata[22:12] == 1833) begin 
      x02bai <= 32'b00111111100001110001001011010101;
      x02jyou <= 32'b00111110100011101000100110111100;
    end else if (wbdata[22:12] == 1834) begin 
      x02bai <= 32'b00111111100001110000100111101101;
      x02jyou <= 32'b00111110100011100111011011110001;
    end else if (wbdata[22:12] == 1835) begin 
      x02bai <= 32'b00111111100001110000000100000110;
      x02jyou <= 32'b00111110100011100110010000101001;
    end else if (wbdata[22:12] == 1836) begin 
      x02bai <= 32'b00111111100001101111100000100000;
      x02jyou <= 32'b00111110100011100101000101100100;
    end else if (wbdata[22:12] == 1837) begin 
      x02bai <= 32'b00111111100001101110111100111100;
      x02jyou <= 32'b00111110100011100011111010100101;
    end else if (wbdata[22:12] == 1838) begin 
      x02bai <= 32'b00111111100001101110011001011000;
      x02jyou <= 32'b00111110100011100010101111100111;
    end else if (wbdata[22:12] == 1839) begin 
      x02bai <= 32'b00111111100001101101110101110110;
      x02jyou <= 32'b00111110100011100001100100101110;
    end else if (wbdata[22:12] == 1840) begin 
      x02bai <= 32'b00111111100001101101010010010101;
      x02jyou <= 32'b00111110100011100000011001111001;
    end else if (wbdata[22:12] == 1841) begin 
      x02bai <= 32'b00111111100001101100101110110101;
      x02jyou <= 32'b00111110100011011111001111000111;
    end else if (wbdata[22:12] == 1842) begin 
      x02bai <= 32'b00111111100001101100001011010111;
      x02jyou <= 32'b00111110100011011110000100011011;
    end else if (wbdata[22:12] == 1843) begin 
      x02bai <= 32'b00111111100001101011100111111001;
      x02jyou <= 32'b00111110100011011100111001110000;
    end else if (wbdata[22:12] == 1844) begin 
      x02bai <= 32'b00111111100001101011000100011101;
      x02jyou <= 32'b00111110100011011011101111001010;
    end else if (wbdata[22:12] == 1845) begin 
      x02bai <= 32'b00111111100001101010100001000010;
      x02jyou <= 32'b00111110100011011010100100100111;
    end else if (wbdata[22:12] == 1846) begin 
      x02bai <= 32'b00111111100001101001111101101000;
      x02jyou <= 32'b00111110100011011001011010001000;
    end else if (wbdata[22:12] == 1847) begin 
      x02bai <= 32'b00111111100001101001011010001111;
      x02jyou <= 32'b00111110100011011000001111101100;
    end else if (wbdata[22:12] == 1848) begin 
      x02bai <= 32'b00111111100001101000110110110111;
      x02jyou <= 32'b00111110100011010111000101010100;
    end else if (wbdata[22:12] == 1849) begin 
      x02bai <= 32'b00111111100001101000010011100001;
      x02jyou <= 32'b00111110100011010101111011000001;
    end else if (wbdata[22:12] == 1850) begin 
      x02bai <= 32'b00111111100001100111110000001011;
      x02jyou <= 32'b00111110100011010100110000101111;
    end else if (wbdata[22:12] == 1851) begin 
      x02bai <= 32'b00111111100001100111001100110111;
      x02jyou <= 32'b00111110100011010011100110100011;
    end else if (wbdata[22:12] == 1852) begin 
      x02bai <= 32'b00111111100001100110101001100100;
      x02jyou <= 32'b00111110100011010010011100011010;
    end else if (wbdata[22:12] == 1853) begin 
      x02bai <= 32'b00111111100001100110000110010010;
      x02jyou <= 32'b00111110100011010001010010010100;
    end else if (wbdata[22:12] == 1854) begin 
      x02bai <= 32'b00111111100001100101100011000010;
      x02jyou <= 32'b00111110100011010000001000010100;
    end else if (wbdata[22:12] == 1855) begin 
      x02bai <= 32'b00111111100001100100111111110010;
      x02jyou <= 32'b00111110100011001110111110010101;
    end else if (wbdata[22:12] == 1856) begin 
      x02bai <= 32'b00111111100001100100011100100100;
      x02jyou <= 32'b00111110100011001101110100011011;
    end else if (wbdata[22:12] == 1857) begin 
      x02bai <= 32'b00111111100001100011111001010110;
      x02jyou <= 32'b00111110100011001100101010100010;
    end else if (wbdata[22:12] == 1858) begin 
      x02bai <= 32'b00111111100001100011010110001010;
      x02jyou <= 32'b00111110100011001011100000101111;
    end else if (wbdata[22:12] == 1859) begin 
      x02bai <= 32'b00111111100001100010110010111111;
      x02jyou <= 32'b00111110100011001010010111000000;
    end else if (wbdata[22:12] == 1860) begin 
      x02bai <= 32'b00111111100001100010001111110110;
      x02jyou <= 32'b00111110100011001001001101010101;
    end else if (wbdata[22:12] == 1861) begin 
      x02bai <= 32'b00111111100001100001101100101101;
      x02jyou <= 32'b00111110100011001000000011101100;
    end else if (wbdata[22:12] == 1862) begin 
      x02bai <= 32'b00111111100001100001001001100101;
      x02jyou <= 32'b00111110100011000110111010000110;
    end else if (wbdata[22:12] == 1863) begin 
      x02bai <= 32'b00111111100001100000100110011111;
      x02jyou <= 32'b00111110100011000101110000100110;
    end else if (wbdata[22:12] == 1864) begin 
      x02bai <= 32'b00111111100001100000000011011010;
      x02jyou <= 32'b00111110100011000100100111001000;
    end else if (wbdata[22:12] == 1865) begin 
      x02bai <= 32'b00111111100001011111100000010110;
      x02jyou <= 32'b00111110100011000011011101101111;
    end else if (wbdata[22:12] == 1866) begin 
      x02bai <= 32'b00111111100001011110111101010011;
      x02jyou <= 32'b00111110100011000010010100011000;
    end else if (wbdata[22:12] == 1867) begin 
      x02bai <= 32'b00111111100001011110011010010001;
      x02jyou <= 32'b00111110100011000001001011000101;
    end else if (wbdata[22:12] == 1868) begin 
      x02bai <= 32'b00111111100001011101110111010001;
      x02jyou <= 32'b00111110100011000000000001110111;
    end else if (wbdata[22:12] == 1869) begin 
      x02bai <= 32'b00111111100001011101010100010001;
      x02jyou <= 32'b00111110100010111110111000101010;
    end else if (wbdata[22:12] == 1870) begin 
      x02bai <= 32'b00111111100001011100110001010011;
      x02jyou <= 32'b00111110100010111101101111100011;
    end else if (wbdata[22:12] == 1871) begin 
      x02bai <= 32'b00111111100001011100001110010110;
      x02jyou <= 32'b00111110100010111100100110011111;
    end else if (wbdata[22:12] == 1872) begin 
      x02bai <= 32'b00111111100001011011101011011010;
      x02jyou <= 32'b00111110100010111011011101011110;
    end else if (wbdata[22:12] == 1873) begin 
      x02bai <= 32'b00111111100001011011001000011111;
      x02jyou <= 32'b00111110100010111010010100100000;
    end else if (wbdata[22:12] == 1874) begin 
      x02bai <= 32'b00111111100001011010100101100101;
      x02jyou <= 32'b00111110100010111001001011100110;
    end else if (wbdata[22:12] == 1875) begin 
      x02bai <= 32'b00111111100001011010000010101100;
      x02jyou <= 32'b00111110100010111000000010101111;
    end else if (wbdata[22:12] == 1876) begin 
      x02bai <= 32'b00111111100001011001011111110101;
      x02jyou <= 32'b00111110100010110110111001111110;
    end else if (wbdata[22:12] == 1877) begin 
      x02bai <= 32'b00111111100001011000111100111111;
      x02jyou <= 32'b00111110100010110101110001001111;
    end else if (wbdata[22:12] == 1878) begin 
      x02bai <= 32'b00111111100001011000011010001001;
      x02jyou <= 32'b00111110100010110100101000100010;
    end else if (wbdata[22:12] == 1879) begin 
      x02bai <= 32'b00111111100001010111110111010101;
      x02jyou <= 32'b00111110100010110011011111111010;
    end else if (wbdata[22:12] == 1880) begin 
      x02bai <= 32'b00111111100001010111010100100010;
      x02jyou <= 32'b00111110100010110010010111010110;
    end else if (wbdata[22:12] == 1881) begin 
      x02bai <= 32'b00111111100001010110110001110001;
      x02jyou <= 32'b00111110100010110001001110110111;
    end else if (wbdata[22:12] == 1882) begin 
      x02bai <= 32'b00111111100001010110001111000000;
      x02jyou <= 32'b00111110100010110000000110011001;
    end else if (wbdata[22:12] == 1883) begin 
      x02bai <= 32'b00111111100001010101101100010000;
      x02jyou <= 32'b00111110100010101110111101111110;
    end else if (wbdata[22:12] == 1884) begin 
      x02bai <= 32'b00111111100001010101001001100010;
      x02jyou <= 32'b00111110100010101101110101101001;
    end else if (wbdata[22:12] == 1885) begin 
      x02bai <= 32'b00111111100001010100100110110101;
      x02jyou <= 32'b00111110100010101100101101010111;
    end else if (wbdata[22:12] == 1886) begin 
      x02bai <= 32'b00111111100001010100000100001001;
      x02jyou <= 32'b00111110100010101011100101001000;
    end else if (wbdata[22:12] == 1887) begin 
      x02bai <= 32'b00111111100001010011100001011110;
      x02jyou <= 32'b00111110100010101010011100111100;
    end else if (wbdata[22:12] == 1888) begin 
      x02bai <= 32'b00111111100001010010111110110100;
      x02jyou <= 32'b00111110100010101001010100110100;
    end else if (wbdata[22:12] == 1889) begin 
      x02bai <= 32'b00111111100001010010011100001011;
      x02jyou <= 32'b00111110100010101000001100101111;
    end else if (wbdata[22:12] == 1890) begin 
      x02bai <= 32'b00111111100001010001111001100011;
      x02jyou <= 32'b00111110100010100111000100101101;
    end else if (wbdata[22:12] == 1891) begin 
      x02bai <= 32'b00111111100001010001010110111101;
      x02jyou <= 32'b00111110100010100101111100110000;
    end else if (wbdata[22:12] == 1892) begin 
      x02bai <= 32'b00111111100001010000110100010111;
      x02jyou <= 32'b00111110100010100100110100110101;
    end else if (wbdata[22:12] == 1893) begin 
      x02bai <= 32'b00111111100001010000010001110011;
      x02jyou <= 32'b00111110100010100011101100111111;
    end else if (wbdata[22:12] == 1894) begin 
      x02bai <= 32'b00111111100001001111101111010000;
      x02jyou <= 32'b00111110100010100010100101001100;
    end else if (wbdata[22:12] == 1895) begin 
      x02bai <= 32'b00111111100001001111001100101110;
      x02jyou <= 32'b00111110100010100001011101011101;
    end else if (wbdata[22:12] == 1896) begin 
      x02bai <= 32'b00111111100001001110101010001101;
      x02jyou <= 32'b00111110100010100000010101110001;
    end else if (wbdata[22:12] == 1897) begin 
      x02bai <= 32'b00111111100001001110000111101101;
      x02jyou <= 32'b00111110100010011111001110001000;
    end else if (wbdata[22:12] == 1898) begin 
      x02bai <= 32'b00111111100001001101100101001111;
      x02jyou <= 32'b00111110100010011110000110100100;
    end else if (wbdata[22:12] == 1899) begin 
      x02bai <= 32'b00111111100001001101000010110001;
      x02jyou <= 32'b00111110100010011100111111000001;
    end else if (wbdata[22:12] == 1900) begin 
      x02bai <= 32'b00111111100001001100100000010101;
      x02jyou <= 32'b00111110100010011011110111100100;
    end else if (wbdata[22:12] == 1901) begin 
      x02bai <= 32'b00111111100001001011111101111001;
      x02jyou <= 32'b00111110100010011010110000001000;
    end else if (wbdata[22:12] == 1902) begin 
      x02bai <= 32'b00111111100001001011011011011111;
      x02jyou <= 32'b00111110100010011001101000110001;
    end else if (wbdata[22:12] == 1903) begin 
      x02bai <= 32'b00111111100001001010111001000110;
      x02jyou <= 32'b00111110100010011000100001011110;
    end else if (wbdata[22:12] == 1904) begin 
      x02bai <= 32'b00111111100001001010010110101110;
      x02jyou <= 32'b00111110100010010111011010001101;
    end else if (wbdata[22:12] == 1905) begin 
      x02bai <= 32'b00111111100001001001110100010111;
      x02jyou <= 32'b00111110100010010110010011000000;
    end else if (wbdata[22:12] == 1906) begin 
      x02bai <= 32'b00111111100001001001010010000001;
      x02jyou <= 32'b00111110100010010101001011110110;
    end else if (wbdata[22:12] == 1907) begin 
      x02bai <= 32'b00111111100001001000101111101101;
      x02jyou <= 32'b00111110100010010100000100110010;
    end else if (wbdata[22:12] == 1908) begin 
      x02bai <= 32'b00111111100001001000001101011001;
      x02jyou <= 32'b00111110100010010010111101101110;
    end else if (wbdata[22:12] == 1909) begin 
      x02bai <= 32'b00111111100001000111101011000111;
      x02jyou <= 32'b00111110100010010001110110110000;
    end else if (wbdata[22:12] == 1910) begin 
      x02bai <= 32'b00111111100001000111001000110110;
      x02jyou <= 32'b00111110100010010000101111110101;
    end else if (wbdata[22:12] == 1911) begin 
      x02bai <= 32'b00111111100001000110100110100101;
      x02jyou <= 32'b00111110100010001111101000111100;
    end else if (wbdata[22:12] == 1912) begin 
      x02bai <= 32'b00111111100001000110000100010110;
      x02jyou <= 32'b00111110100010001110100010000111;
    end else if (wbdata[22:12] == 1913) begin 
      x02bai <= 32'b00111111100001000101100010001000;
      x02jyou <= 32'b00111110100010001101011011010110;
    end else if (wbdata[22:12] == 1914) begin 
      x02bai <= 32'b00111111100001000100111111111011;
      x02jyou <= 32'b00111110100010001100010100101000;
    end else if (wbdata[22:12] == 1915) begin 
      x02bai <= 32'b00111111100001000100011101110000;
      x02jyou <= 32'b00111110100010001011001101111111;
    end else if (wbdata[22:12] == 1916) begin 
      x02bai <= 32'b00111111100001000011111011100101;
      x02jyou <= 32'b00111110100010001010000111010111;
    end else if (wbdata[22:12] == 1917) begin 
      x02bai <= 32'b00111111100001000011011001011011;
      x02jyou <= 32'b00111110100010001001000000110011;
    end else if (wbdata[22:12] == 1918) begin 
      x02bai <= 32'b00111111100001000010110111010011;
      x02jyou <= 32'b00111110100010000111111010010100;
    end else if (wbdata[22:12] == 1919) begin 
      x02bai <= 32'b00111111100001000010010101001100;
      x02jyou <= 32'b00111110100010000110110011111000;
    end else if (wbdata[22:12] == 1920) begin 
      x02bai <= 32'b00111111100001000001110011000101;
      x02jyou <= 32'b00111110100010000101101101011101;
    end else if (wbdata[22:12] == 1921) begin 
      x02bai <= 32'b00111111100001000001010001000000;
      x02jyou <= 32'b00111110100010000100100111000111;
    end else if (wbdata[22:12] == 1922) begin 
      x02bai <= 32'b00111111100001000000101110111100;
      x02jyou <= 32'b00111110100010000011100000110101;
    end else if (wbdata[22:12] == 1923) begin 
      x02bai <= 32'b00111111100001000000001100111001;
      x02jyou <= 32'b00111110100010000010011010100110;
    end else if (wbdata[22:12] == 1924) begin 
      x02bai <= 32'b00111111100000111111101010110111;
      x02jyou <= 32'b00111110100010000001010100011010;
    end else if (wbdata[22:12] == 1925) begin 
      x02bai <= 32'b00111111100000111111001000110111;
      x02jyou <= 32'b00111110100010000000001110010011;
    end else if (wbdata[22:12] == 1926) begin 
      x02bai <= 32'b00111111100000111110100110110111;
      x02jyou <= 32'b00111110100001111111001000001101;
    end else if (wbdata[22:12] == 1927) begin 
      x02bai <= 32'b00111111100000111110000100111000;
      x02jyou <= 32'b00111110100001111110000010001011;
    end else if (wbdata[22:12] == 1928) begin 
      x02bai <= 32'b00111111100000111101100010111011;
      x02jyou <= 32'b00111110100001111100111100001110;
    end else if (wbdata[22:12] == 1929) begin 
      x02bai <= 32'b00111111100000111101000000111110;
      x02jyou <= 32'b00111110100001111011110110010010;
    end else if (wbdata[22:12] == 1930) begin 
      x02bai <= 32'b00111111100000111100011111000011;
      x02jyou <= 32'b00111110100001111010110000011011;
    end else if (wbdata[22:12] == 1931) begin 
      x02bai <= 32'b00111111100000111011111101001001;
      x02jyou <= 32'b00111110100001111001101010100111;
    end else if (wbdata[22:12] == 1932) begin 
      x02bai <= 32'b00111111100000111011011011010000;
      x02jyou <= 32'b00111110100001111000100100110111;
    end else if (wbdata[22:12] == 1933) begin 
      x02bai <= 32'b00111111100000111010111001011000;
      x02jyou <= 32'b00111110100001110111011111001010;
    end else if (wbdata[22:12] == 1934) begin 
      x02bai <= 32'b00111111100000111010010111100001;
      x02jyou <= 32'b00111110100001110110011001100000;
    end else if (wbdata[22:12] == 1935) begin 
      x02bai <= 32'b00111111100000111001110101101011;
      x02jyou <= 32'b00111110100001110101010011111001;
    end else if (wbdata[22:12] == 1936) begin 
      x02bai <= 32'b00111111100000111001010011110110;
      x02jyou <= 32'b00111110100001110100001110010101;
    end else if (wbdata[22:12] == 1937) begin 
      x02bai <= 32'b00111111100000111000110010000011;
      x02jyou <= 32'b00111110100001110011001000110110;
    end else if (wbdata[22:12] == 1938) begin 
      x02bai <= 32'b00111111100000111000010000010000;
      x02jyou <= 32'b00111110100001110010000011011001;
    end else if (wbdata[22:12] == 1939) begin 
      x02bai <= 32'b00111111100000110111101110011110;
      x02jyou <= 32'b00111110100001110000111101111111;
    end else if (wbdata[22:12] == 1940) begin 
      x02bai <= 32'b00111111100000110111001100101110;
      x02jyou <= 32'b00111110100001101111111000101010;
    end else if (wbdata[22:12] == 1941) begin 
      x02bai <= 32'b00111111100000110110101010111111;
      x02jyou <= 32'b00111110100001101110110011011000;
    end else if (wbdata[22:12] == 1942) begin 
      x02bai <= 32'b00111111100000110110001001010000;
      x02jyou <= 32'b00111110100001101101101110000111;
    end else if (wbdata[22:12] == 1943) begin 
      x02bai <= 32'b00111111100000110101100111100011;
      x02jyou <= 32'b00111110100001101100101000111100;
    end else if (wbdata[22:12] == 1944) begin 
      x02bai <= 32'b00111111100000110101000101110111;
      x02jyou <= 32'b00111110100001101011100011110011;
    end else if (wbdata[22:12] == 1945) begin 
      x02bai <= 32'b00111111100000110100100100001100;
      x02jyou <= 32'b00111110100001101010011110101110;
    end else if (wbdata[22:12] == 1946) begin 
      x02bai <= 32'b00111111100000110100000010100010;
      x02jyou <= 32'b00111110100001101001011001101100;
    end else if (wbdata[22:12] == 1947) begin 
      x02bai <= 32'b00111111100000110011100000111001;
      x02jyou <= 32'b00111110100001101000010100101101;
    end else if (wbdata[22:12] == 1948) begin 
      x02bai <= 32'b00111111100000110010111111010010;
      x02jyou <= 32'b00111110100001100111001111110100;
    end else if (wbdata[22:12] == 1949) begin 
      x02bai <= 32'b00111111100000110010011101101011;
      x02jyou <= 32'b00111110100001100110001010111011;
    end else if (wbdata[22:12] == 1950) begin 
      x02bai <= 32'b00111111100000110001111100000101;
      x02jyou <= 32'b00111110100001100101000110000110;
    end else if (wbdata[22:12] == 1951) begin 
      x02bai <= 32'b00111111100000110001011010100001;
      x02jyou <= 32'b00111110100001100100000001010110;
    end else if (wbdata[22:12] == 1952) begin 
      x02bai <= 32'b00111111100000110000111000111101;
      x02jyou <= 32'b00111110100001100010111100100110;
    end else if (wbdata[22:12] == 1953) begin 
      x02bai <= 32'b00111111100000110000010111011011;
      x02jyou <= 32'b00111110100001100001110111111101;
    end else if (wbdata[22:12] == 1954) begin 
      x02bai <= 32'b00111111100000101111110101111001;
      x02jyou <= 32'b00111110100001100000110011010100;
    end else if (wbdata[22:12] == 1955) begin 
      x02bai <= 32'b00111111100000101111010100011001;
      x02jyou <= 32'b00111110100001011111101110110000;
    end else if (wbdata[22:12] == 1956) begin 
      x02bai <= 32'b00111111100000101110110010111010;
      x02jyou <= 32'b00111110100001011110101010010000;
    end else if (wbdata[22:12] == 1957) begin 
      x02bai <= 32'b00111111100000101110010001011100;
      x02jyou <= 32'b00111110100001011101100101110010;
    end else if (wbdata[22:12] == 1958) begin 
      x02bai <= 32'b00111111100000101101101111111111;
      x02jyou <= 32'b00111110100001011100100001011000;
    end else if (wbdata[22:12] == 1959) begin 
      x02bai <= 32'b00111111100000101101001110100011;
      x02jyou <= 32'b00111110100001011011011101000001;
    end else if (wbdata[22:12] == 1960) begin 
      x02bai <= 32'b00111111100000101100101101001000;
      x02jyou <= 32'b00111110100001011010011000101101;
    end else if (wbdata[22:12] == 1961) begin 
      x02bai <= 32'b00111111100000101100001011101110;
      x02jyou <= 32'b00111110100001011001010100011100;
    end else if (wbdata[22:12] == 1962) begin 
      x02bai <= 32'b00111111100000101011101010010101;
      x02jyou <= 32'b00111110100001011000010000001111;
    end else if (wbdata[22:12] == 1963) begin 
      x02bai <= 32'b00111111100000101011001000111101;
      x02jyou <= 32'b00111110100001010111001100000100;
    end else if (wbdata[22:12] == 1964) begin 
      x02bai <= 32'b00111111100000101010100111100111;
      x02jyou <= 32'b00111110100001010110000111111111;
    end else if (wbdata[22:12] == 1965) begin 
      x02bai <= 32'b00111111100000101010000110010001;
      x02jyou <= 32'b00111110100001010101000011111010;
    end else if (wbdata[22:12] == 1966) begin 
      x02bai <= 32'b00111111100000101001100100111101;
      x02jyou <= 32'b00111110100001010011111111111011;
    end else if (wbdata[22:12] == 1967) begin 
      x02bai <= 32'b00111111100000101001000011101001;
      x02jyou <= 32'b00111110100001010010111011111101;
    end else if (wbdata[22:12] == 1968) begin 
      x02bai <= 32'b00111111100000101000100010010111;
      x02jyou <= 32'b00111110100001010001111000000100;
    end else if (wbdata[22:12] == 1969) begin 
      x02bai <= 32'b00111111100000101000000001000101;
      x02jyou <= 32'b00111110100001010000110100001101;
    end else if (wbdata[22:12] == 1970) begin 
      x02bai <= 32'b00111111100000100111011111110101;
      x02jyou <= 32'b00111110100001001111110000011010;
    end else if (wbdata[22:12] == 1971) begin 
      x02bai <= 32'b00111111100000100110111110100110;
      x02jyou <= 32'b00111110100001001110101100101011;
    end else if (wbdata[22:12] == 1972) begin 
      x02bai <= 32'b00111111100000100110011101011000;
      x02jyou <= 32'b00111110100001001101101000111110;
    end else if (wbdata[22:12] == 1973) begin 
      x02bai <= 32'b00111111100000100101111100001011;
      x02jyou <= 32'b00111110100001001100100101010101;
    end else if (wbdata[22:12] == 1974) begin 
      x02bai <= 32'b00111111100000100101011010111111;
      x02jyou <= 32'b00111110100001001011100001101111;
    end else if (wbdata[22:12] == 1975) begin 
      x02bai <= 32'b00111111100000100100111001110100;
      x02jyou <= 32'b00111110100001001010011110001100;
    end else if (wbdata[22:12] == 1976) begin 
      x02bai <= 32'b00111111100000100100011000101010;
      x02jyou <= 32'b00111110100001001001011010101100;
    end else if (wbdata[22:12] == 1977) begin 
      x02bai <= 32'b00111111100000100011110111100001;
      x02jyou <= 32'b00111110100001001000010111001111;
    end else if (wbdata[22:12] == 1978) begin 
      x02bai <= 32'b00111111100000100011010110011001;
      x02jyou <= 32'b00111110100001000111010011110101;
    end else if (wbdata[22:12] == 1979) begin 
      x02bai <= 32'b00111111100000100010110101010010;
      x02jyou <= 32'b00111110100001000110010000011111;
    end else if (wbdata[22:12] == 1980) begin 
      x02bai <= 32'b00111111100000100010010100001100;
      x02jyou <= 32'b00111110100001000101001101001011;
    end else if (wbdata[22:12] == 1981) begin 
      x02bai <= 32'b00111111100000100001110011001000;
      x02jyou <= 32'b00111110100001000100001001111101;
    end else if (wbdata[22:12] == 1982) begin 
      x02bai <= 32'b00111111100000100001010010000100;
      x02jyou <= 32'b00111110100001000011000110101111;
    end else if (wbdata[22:12] == 1983) begin 
      x02bai <= 32'b00111111100000100000110001000010;
      x02jyou <= 32'b00111110100001000010000011100111;
    end else if (wbdata[22:12] == 1984) begin 
      x02bai <= 32'b00111111100000100000010000000000;
      x02jyou <= 32'b00111110100001000001000000100000;
    end else if (wbdata[22:12] == 1985) begin 
      x02bai <= 32'b00111111100000011111101111000000;
      x02jyou <= 32'b00111110100000111111111101011110;
    end else if (wbdata[22:12] == 1986) begin 
      x02bai <= 32'b00111111100000011111001110000000;
      x02jyou <= 32'b00111110100000111110111010011101;
    end else if (wbdata[22:12] == 1987) begin 
      x02bai <= 32'b00111111100000011110101101000010;
      x02jyou <= 32'b00111110100000111101110111100001;
    end else if (wbdata[22:12] == 1988) begin 
      x02bai <= 32'b00111111100000011110001100000100;
      x02jyou <= 32'b00111110100000111100110100100111;
    end else if (wbdata[22:12] == 1989) begin 
      x02bai <= 32'b00111111100000011101101011001000;
      x02jyou <= 32'b00111110100000111011110001110001;
    end else if (wbdata[22:12] == 1990) begin 
      x02bai <= 32'b00111111100000011101001010001101;
      x02jyou <= 32'b00111110100000111010101110111111;
    end else if (wbdata[22:12] == 1991) begin 
      x02bai <= 32'b00111111100000011100101001010011;
      x02jyou <= 32'b00111110100000111001101100001111;
    end else if (wbdata[22:12] == 1992) begin 
      x02bai <= 32'b00111111100000011100001000011001;
      x02jyou <= 32'b00111110100000111000101001100001;
    end else if (wbdata[22:12] == 1993) begin 
      x02bai <= 32'b00111111100000011011100111100001;
      x02jyou <= 32'b00111110100000110111100110110111;
    end else if (wbdata[22:12] == 1994) begin 
      x02bai <= 32'b00111111100000011011000110101010;
      x02jyou <= 32'b00111110100000110110100100010001;
    end else if (wbdata[22:12] == 1995) begin 
      x02bai <= 32'b00111111100000011010100101110100;
      x02jyou <= 32'b00111110100000110101100001101110;
    end else if (wbdata[22:12] == 1996) begin 
      x02bai <= 32'b00111111100000011010000100111111;
      x02jyou <= 32'b00111110100000110100011111001110;
    end else if (wbdata[22:12] == 1997) begin 
      x02bai <= 32'b00111111100000011001100100001011;
      x02jyou <= 32'b00111110100000110011011100110001;
    end else if (wbdata[22:12] == 1998) begin 
      x02bai <= 32'b00111111100000011001000011011000;
      x02jyou <= 32'b00111110100000110010011010010111;
    end else if (wbdata[22:12] == 1999) begin 
      x02bai <= 32'b00111111100000011000100010100110;
      x02jyou <= 32'b00111110100000110001011000000000;
    end else if (wbdata[22:12] == 2000) begin 
      x02bai <= 32'b00111111100000011000000001110101;
      x02jyou <= 32'b00111110100000110000010101101101;
    end else if (wbdata[22:12] == 2001) begin 
      x02bai <= 32'b00111111100000010111100001000110;
      x02jyou <= 32'b00111110100000101111010011011110;
    end else if (wbdata[22:12] == 2002) begin 
      x02bai <= 32'b00111111100000010111000000010111;
      x02jyou <= 32'b00111110100000101110010001010001;
    end else if (wbdata[22:12] == 2003) begin 
      x02bai <= 32'b00111111100000010110011111101001;
      x02jyou <= 32'b00111110100000101101001111000110;
    end else if (wbdata[22:12] == 2004) begin 
      x02bai <= 32'b00111111100000010101111110111100;
      x02jyou <= 32'b00111110100000101100001100111111;
    end else if (wbdata[22:12] == 2005) begin 
      x02bai <= 32'b00111111100000010101011110010001;
      x02jyou <= 32'b00111110100000101011001010111100;
    end else if (wbdata[22:12] == 2006) begin 
      x02bai <= 32'b00111111100000010100111101100110;
      x02jyou <= 32'b00111110100000101010001000111011;
    end else if (wbdata[22:12] == 2007) begin 
      x02bai <= 32'b00111111100000010100011100111100;
      x02jyou <= 32'b00111110100000101001000110111101;
    end else if (wbdata[22:12] == 2008) begin 
      x02bai <= 32'b00111111100000010011111100010100;
      x02jyou <= 32'b00111110100000101000000101000011;
    end else if (wbdata[22:12] == 2009) begin 
      x02bai <= 32'b00111111100000010011011011101100;
      x02jyou <= 32'b00111110100000100111000011001011;
    end else if (wbdata[22:12] == 2010) begin 
      x02bai <= 32'b00111111100000010010111011000110;
      x02jyou <= 32'b00111110100000100110000001011000;
    end else if (wbdata[22:12] == 2011) begin 
      x02bai <= 32'b00111111100000010010011010100000;
      x02jyou <= 32'b00111110100000100100111111100110;
    end else if (wbdata[22:12] == 2012) begin 
      x02bai <= 32'b00111111100000010001111001111100;
      x02jyou <= 32'b00111110100000100011111101111001;
    end else if (wbdata[22:12] == 2013) begin 
      x02bai <= 32'b00111111100000010001011001011000;
      x02jyou <= 32'b00111110100000100010111100001101;
    end else if (wbdata[22:12] == 2014) begin 
      x02bai <= 32'b00111111100000010000111000110110;
      x02jyou <= 32'b00111110100000100001111010100110;
    end else if (wbdata[22:12] == 2015) begin 
      x02bai <= 32'b00111111100000010000011000010100;
      x02jyou <= 32'b00111110100000100000111001000001;
    end else if (wbdata[22:12] == 2016) begin 
      x02bai <= 32'b00111111100000001111110111110100;
      x02jyou <= 32'b00111110100000011111110111100000;
    end else if (wbdata[22:12] == 2017) begin 
      x02bai <= 32'b00111111100000001111010111010101;
      x02jyou <= 32'b00111110100000011110110110000010;
    end else if (wbdata[22:12] == 2018) begin 
      x02bai <= 32'b00111111100000001110110110110110;
      x02jyou <= 32'b00111110100000011101110100100101;
    end else if (wbdata[22:12] == 2019) begin 
      x02bai <= 32'b00111111100000001110010110011001;
      x02jyou <= 32'b00111110100000011100110011001110;
    end else if (wbdata[22:12] == 2020) begin 
      x02bai <= 32'b00111111100000001101110101111101;
      x02jyou <= 32'b00111110100000011011110001111001;
    end else if (wbdata[22:12] == 2021) begin 
      x02bai <= 32'b00111111100000001101010101100010;
      x02jyou <= 32'b00111110100000011010110000101000;
    end else if (wbdata[22:12] == 2022) begin 
      x02bai <= 32'b00111111100000001100110101000111;
      x02jyou <= 32'b00111110100000011001101111010111;
    end else if (wbdata[22:12] == 2023) begin 
      x02bai <= 32'b00111111100000001100010100101110;
      x02jyou <= 32'b00111110100000011000101110001100;
    end else if (wbdata[22:12] == 2024) begin 
      x02bai <= 32'b00111111100000001011110100010110;
      x02jyou <= 32'b00111110100000010111101101000011;
    end else if (wbdata[22:12] == 2025) begin 
      x02bai <= 32'b00111111100000001011010011111111;
      x02jyou <= 32'b00111110100000010110101011111110;
    end else if (wbdata[22:12] == 2026) begin 
      x02bai <= 32'b00111111100000001010110011101000;
      x02jyou <= 32'b00111110100000010101101010111010;
    end else if (wbdata[22:12] == 2027) begin 
      x02bai <= 32'b00111111100000001010010011010011;
      x02jyou <= 32'b00111110100000010100101001111010;
    end else if (wbdata[22:12] == 2028) begin 
      x02bai <= 32'b00111111100000001001110010111111;
      x02jyou <= 32'b00111110100000010011101000111110;
    end else if (wbdata[22:12] == 2029) begin 
      x02bai <= 32'b00111111100000001001010010101100;
      x02jyou <= 32'b00111110100000010010101000000101;
    end else if (wbdata[22:12] == 2030) begin 
      x02bai <= 32'b00111111100000001000110010011010;
      x02jyou <= 32'b00111110100000010001100111001110;
    end else if (wbdata[22:12] == 2031) begin 
      x02bai <= 32'b00111111100000001000010010001001;
      x02jyou <= 32'b00111110100000010000100110011011;
    end else if (wbdata[22:12] == 2032) begin 
      x02bai <= 32'b00111111100000000111110001111001;
      x02jyou <= 32'b00111110100000001111100101101011;
    end else if (wbdata[22:12] == 2033) begin 
      x02bai <= 32'b00111111100000000111010001101010;
      x02jyou <= 32'b00111110100000001110100100111110;
    end else if (wbdata[22:12] == 2034) begin 
      x02bai <= 32'b00111111100000000110110001011100;
      x02jyou <= 32'b00111110100000001101100100010100;
    end else if (wbdata[22:12] == 2035) begin 
      x02bai <= 32'b00111111100000000110010001001110;
      x02jyou <= 32'b00111110100000001100100011101011;
    end else if (wbdata[22:12] == 2036) begin 
      x02bai <= 32'b00111111100000000101110001000010;
      x02jyou <= 32'b00111110100000001011100011000110;
    end else if (wbdata[22:12] == 2037) begin 
      x02bai <= 32'b00111111100000000101010000110111;
      x02jyou <= 32'b00111110100000001010100010100101;
    end else if (wbdata[22:12] == 2038) begin 
      x02bai <= 32'b00111111100000000100110000101101;
      x02jyou <= 32'b00111110100000001001100010000111;
    end else if (wbdata[22:12] == 2039) begin 
      x02bai <= 32'b00111111100000000100010000100100;
      x02jyou <= 32'b00111110100000001000100001101100;
    end else if (wbdata[22:12] == 2040) begin 
      x02bai <= 32'b00111111100000000011110000011100;
      x02jyou <= 32'b00111110100000000111100001010100;
    end else if (wbdata[22:12] == 2041) begin 
      x02bai <= 32'b00111111100000000011010000010101;
      x02jyou <= 32'b00111110100000000110100000111111;
    end else if (wbdata[22:12] == 2042) begin 
      x02bai <= 32'b00111111100000000010110000001111;
      x02jyou <= 32'b00111110100000000101100000101101;
    end else if (wbdata[22:12] == 2043) begin 
      x02bai <= 32'b00111111100000000010010000001010;
      x02jyou <= 32'b00111110100000000100100000011110;
    end else if (wbdata[22:12] == 2044) begin 
      x02bai <= 32'b00111111100000000001110000000110;
      x02jyou <= 32'b00111110100000000011100000010010;
    end else if (wbdata[22:12] == 2045) begin 
      x02bai <= 32'b00111111100000000001010000000011;
      x02jyou <= 32'b00111110100000000010100000001001;
    end else if (wbdata[22:12] == 2046) begin 
      x02bai <= 32'b00111111100000000000110000000001;
      x02jyou <= 32'b00111110100000000001100000000011;
    end else if (wbdata[22:12] == 2047) begin 
      x02bai <= 32'b00111111100000000000010000000000;
      x02jyou <= 32'b00111110100000000000100000000000;
    end
  end else if (state == STAGE2) begin
    state <= STAGE3;
    adata2 <= adata1;
    bdata2 <= bdata1;
    x02bai2 <= x02bai;
      ax02s1 <= 1'b0;
      ax02e1 <= 9'd127 + x02jyou[30:23];
      bdatakari <= {1'b1,bdata1[22:0]};
      x2jyoukari <= {1'b1,x02jyou[22:0]};
  end else if (state == STAGE3) begin
    state <= STAGE4;
    adata3 <= adata2;
    bdata3 <= bdata2;
    x02bai3 <= x02bai2;
    ax02jyous2 <= ax02s1;
    ax02jyoue2 <= ax02e1 - 9'd127;
    ax02jyoukekka <= bdatakari * x2jyoukari;
  end else if (state == STAGE4) begin
    state <= STAGE5;
    adata4 <= adata3;
    bdata4 <= bdata3;
    x02bai4 <= x02bai3;
    if (ax02jyoukekka[47] == 1) begin
      minusax02jyou <= {~ax02jyous2,ax02jyoue2[7:0]+8'd1,ax02jyoukekka[46:24]};
    end else begin
      minusax02jyou <= {~ax02jyous2,ax02jyoue2[7:0],ax02jyoukekka[45:23]};
    end
  end else if (state == STAGE5) begin
        state <= STAGE6;
        adata5 <= adata4;
        bdata5 <= bdata4;
    if (x02bai4[31] == minusax02jyou[31]) begin
      invbtashi1hiki0 <= 1;
    end else begin
      invbtashi1hiki0 <= 0;
    end
    if ((x02bai4[30:23] > minusax02jyou[30:23]) || ((x02bai4[30:23] == minusax02jyou[30:23]) && (x02bai4[22:0] >= minusax02jyou[22:0]))) begin
      invbs1 <= x02bai4[31];
      invbe1 <= x02bai4[30:23];
      invbdeka <= {1'b0,1'b1,x02bai4[22:0]};
      invbchibi <= ({1'b0,1'b1,minusax02jyou[22:0]} >> (x02bai4[30:23] - minusax02jyou[30:23]));
    end else begin
      invbs1 <= minusax02jyou[31];
      invbe1 <= minusax02jyou[30:23];
      invbdeka <= {1'b0,1'b1,minusax02jyou[22:0]};
      invbchibi <= ({1'b0,1'b1,x02bai4[22:0]} >> (minusax02jyou[30:23] - x02bai4[30:23]));
    end
  end else if (state == STAGE6) begin
    state <= STAGE7;
    adata6 <= adata5;
    bdata6 <= bdata5;
    invbs2 <= invbs1;
    invbe2 <= invbe1;
    if (invbtashi1hiki0 == 1) begin
      invbkekka <= invbdeka[24:0] + invbchibi[24:0];
    end else begin
      invbkekka <= invbdeka[24:0] - invbchibi[24:0];
    end
  end else if (state == STAGE7) begin
    state <= STAGE8;
    adata7 <= adata6;
    bdata7 <= bdata6;
    if (invbkekka[24] == 1) begin
      invb <= {invbs2,invbe2[7:0]+8'd1,invbkekka[23:1]};
    end else if (invbkekka[23] == 1) begin
      invb <= {invbs2,invbe2[7:0],invbkekka[22:0]};
    end else if (invbkekka[22] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd1,invbkekka[21:0],1'b0};
    end else if (invbkekka[21] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd2,invbkekka[20:0],2'b0};
    end else if (invbkekka[20] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd3,invbkekka[19:0],3'b0};
    end else if (invbkekka[19] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd4,invbkekka[18:0],4'b0};
    end else if (invbkekka[18] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd5,invbkekka[17:0],5'b0};
    end else if (invbkekka[17] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd6,invbkekka[16:0],6'b0};
    end else if (invbkekka[16] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd7,invbkekka[15:0],7'b0};
    end else if (invbkekka[15] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd8,invbkekka[14:0],8'b0};
    end else if (invbkekka[14] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd9,invbkekka[13:0],9'b0};
    end else if (invbkekka[13] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd10,invbkekka[12:0],10'b0};
    end else if (invbkekka[12] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd11,invbkekka[11:0],11'b0};
    end else if (invbkekka[11] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd12,invbkekka[10:0],12'b0};
    end else if (invbkekka[10] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd13,invbkekka[9:0],13'b0};
    end else if (invbkekka[9] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd14,invbkekka[8:0],14'b0};
    end else if (invbkekka[8] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd15,invbkekka[7:0],15'b0};
    end else if (invbkekka[7] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd16,invbkekka[6:0],16'b0};
    end else if (invbkekka[6] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd17,invbkekka[5:0],17'b0};
    end else if (invbkekka[5] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd18,invbkekka[4:0],18'b0};
    end else if (invbkekka[4] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd19,invbkekka[3:0],19'b0};
    end else if (invbkekka[3] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd20,invbkekka[2:0],20'b0};
    end else if (invbkekka[2] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd21,invbkekka[1:0],21'b0};
    end else if (invbkekka[1] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd22,invbkekka[0:0],22'b0};
    end else if (invbkekka[0] == 1) begin
      invb <= {invbs2,invbe2[7:0]-8'd23,23'b0};
    end else begin
      invb <= 0;
    end
  end else if (state == STAGE8) begin
        state <= STAGE9;
      s1 <= adata7[31] ^ bdata7[31];
      e1 <= adata7[30:23] + 9'd127 + invb[30:23];
      esyuuseib <= bdata[30:23];
      if (adata7[30:23] == 0) begin
      if (adata7[22] == 1) begin
	esyuuseia <= 0;
	adatakari <= {adata7[22:0],1'b0};
      end else if (adata7[21] == 1) begin
	esyuuseia <= 1;
	adatakari <= {adata7[21:0],2'b0};
      end else if (adata7[20] == 1) begin
	esyuuseia <= 2;
	adatakari <= {adata7[20:0],3'b0};
      end else if (adata7[19] == 1) begin
	esyuuseia <= 3;
	adatakari <= {adata7[19:0],4'b0};
      end else if (adata7[18] == 1) begin
	esyuuseia <= 4;
	adatakari <= {adata7[18:0],5'b0};
      end else if (adata7[17] == 1) begin
	esyuuseia <= 5;
	adatakari <= {adata7[17:0],6'b0};
      end else if (adata7[16] == 1) begin
	esyuuseia <= 6;
	adatakari <= {adata7[16:0],7'b0};
      end else if (adata7[15] == 1) begin
	esyuuseia <= 7;
	adatakari <= {adata7[15:0],8'b0};
      end else if (adata7[14] == 1) begin
	esyuuseia <= 8;
	adatakari <= {adata7[14:0],9'b0};
      end else if (adata7[13] == 1) begin
	esyuuseia <= 9;
	adatakari <= {adata7[13:0],10'b0};
      end else if (adata7[12] == 1) begin
	esyuuseia <= 10;
	adatakari <= {adata7[12:0],11'b0};
      end else if (adata7[11] == 1) begin
	esyuuseia <= 11;
	adatakari <= {adata7[11:0],12'b0};
      end else if (adata7[10] == 1) begin
	esyuuseia <= 12;
	adatakari <= {adata7[10:0],13'b0};
      end else if (adata7[9] == 1) begin
	esyuuseia <= 13;
	adatakari <= {adata7[9:0],14'b0};
      end else if (adata7[8] == 1) begin
	esyuuseia <= 14;
	adatakari <= {adata7[8:0],15'b0};
      end else if (adata7[7] == 1) begin
	esyuuseia <= 15;
	adatakari <= {adata7[7:0],16'b0};
      end else if (adata7[6] == 1) begin
	esyuuseia <= 16;
	adatakari <= {adata7[6:0],17'b0};
      end else if (adata7[5] == 1) begin
	esyuuseia <= 17;
	adatakari <= {adata7[5:0],18'b0};
      end else if (adata7[4] == 1) begin
	esyuuseia <= 18;
	adatakari <= {adata7[4:0],19'b0};
      end else if (adata7[3] == 1) begin
	esyuuseia <= 19;
	adatakari <= {adata7[3:0],20'b0};
      end else if (adata7[2] == 1) begin
	esyuuseia <= 20;
	adatakari <= {adata7[2:0],21'b0};
      end else if (adata7[1] == 1) begin
	esyuuseia <= 21;
	adatakari <= {adata7[1:0],22'b0};
      end else if (adata7[0] == 1) begin
	esyuuseia <= 22;
	adatakari <= {1'b1,23'b0};
      end else begin
	esyuuseia <= 23;
	adatakari <= 0;
      end
    end else begin
      esyuuseia <= 0;
      adatakari <= {1'b1,adata7[22:0]};
    end
      invbkari <= {1'b1,invb[22:0]};
  end else if (state == STAGE9) begin
    state <= STAGE10;
    s2 <= s1;
    underflow <= (esyuuseia == 23 || (e1 < (esyuuseib + esyuuseia + 127))) ? 1 : 0;
    e2 <=  e1 - esyuuseia - esyuuseib - 9'd127;
    kekka <= adatakari * invbkari;
  end else if (state == STAGE10) begin
    done <= 1;
    busy <= 0;
    state <= WAIT_ST;
    if (underflow == 1) begin
    result <= 32'b0;
    end else
    if (kekka[47] == 1) begin
      result <= {s2,e2[7:0]+8'd1,kekka[46:24]};
    end else begin
      result <= (e2 == 0) ? {s2,8'b0,kekka[46:24]} : {s2,e2[7:0],kekka[45:23]};
    end
  end
end
endmodule

`default_nettype wire


